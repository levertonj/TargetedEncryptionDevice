// crypto_test_tb.v

// Generated using ACDS version 14.1 190 at 2015.03.23.23:35:01

`timescale 1 ps / 1 ps
module crypto_test_tb (
	);

	wire    crypto_test_inst_clk_bfm_clk_clk;       // crypto_test_inst_clk_bfm:clk -> [crypto_test_inst:clk_clk, crypto_test_inst_reset_bfm:clk]
	wire    crypto_test_inst_reset_bfm_reset_reset; // crypto_test_inst_reset_bfm:reset -> crypto_test_inst:reset_reset_n

	crypto_test crypto_test_inst (
		.clk_clk       (crypto_test_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (crypto_test_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) crypto_test_inst_clk_bfm (
		.clk (crypto_test_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) crypto_test_inst_reset_bfm (
		.reset (crypto_test_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (crypto_test_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
