// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
jRtYfiPujijnkEdW25a236eOyOaoCtWlzDgdYET3ucdB32dcMRv9XhKK9Y4wzBiLDl0muga4yP/L
tswXo0SZpNZVetiK5DuSSsMmvmNC+uyKx19k88A3BZ56S+mSY9P7fKb35P9KKiTdPjRfyW9FrAAs
6hcm/CdgScAr2e7yfxXMBWlSnSth6d7FdgZifghlzymOZt7VlA9Cj9BLrQLHfXv+got+DjhNg9Ry
URBussly9BydO80oj5/JS19MmvCZFYkplpHEIR65MopdmwB6LCQnl59xJ8wJGyR4rK92nWSgXtaE
i1ijgc7VoO+ced+JYRJ8jh+RZZVd+kH6ytVhiw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
FFkBoLS+ttgMlXURwur3C7g4CgJV5NQ/q9q/lMPFDqMYXsxq6JX9wpDUxYrAtkgC4FWv63Cgkix3
vQv5hkeN2kuPjhMZZn7wxHmuDGBU+Bn/AvfYujPZ8SLzr4qKlOaDOEaRDyGCDFWtvGcXr20R4iW1
Be8NCUQY0lxWBmruZbnvAePb2psFCXARXFYo0QvO+W0Cj+NJARjFY1NP9mpnujw9EGo4Zg+y/iSu
hjVBxg0UxIRJl8YB2mlE1Vn3+A+Y6Fu2dpmO6VSJBCfjVxbdACnKoMZFcas5piNpmPEp+ZuyxDd/
iFNfik355E2vhwWgg/RbitZ6Pzsv9/rXYkK23MsF8JP6NuSI1e8F9xtH6EKnjKgmfEbUK/rNsdaD
03sk9il24NhHUjvvi5Y7d9nB4mJAiNrChuRExJcgHtCrD1aD1cjGV2dkypPWtQKFlyQuAVjgz2qp
gMcYziv7YYgA4NhZ2VKSaCL4zM3Ghg6RA9OGgByc255FSs9EY62bLnFxJoAxHiGziIaGWWnRYaTj
SupPQt79ZmZZpvZJ8uluCbG6l26+ItZZy/xzcsQlvfCn4zVjDcwjg0lVjsltauMZe6WiE35bZaN7
Yx41Zf+CLk8ZXyAZCjYbVaEdx2W2gAMVlgNTUsZrIeVVBPorPpwQp4lWC77I5tCDjvjzqeNpgoST
f8ws8nEcqXQUQ5uTLaM9dLgnDx4nodwlkgpBwm0d9kj0iU/kOAWH5KJ3jeh3IL2FyL7Y3yGsQKxB
GsMA9PCDyQDUHtop3tRY5UyI1IKyVL58w96bryeNfi9nrpNKWYPPByV4jDKxEWAmjusTMuamjsgf
sBBsSoDfOfUm6lYqzKPApor+dl3r2wCppSxQdPpunUzRBVmVsV2rdZ/1Whvl/aW4QegkQX5HhiZQ
MoCbu7VM6g5ATzPBAtmr5jbpDTjGnxHkdgutnECV3Yc3DlIXwEwZOLPV+6KjoTI2rVzPRq5RRxoz
MKmNeUMazeBsrITb3W0lEiKOGUDKxZyT1LS+qagHsSMWUZykk02iKIyh3LPou4kr/VHV9yac5Tc7
HNwO8Sda37p2JsCBLaat8r0Fdkz/j64UP/re7Ti4tRWPjDQxh+RUEtzfD5t75HwFjX9S7v4/HD5C
zXgGue3kSgfqQ3e+LTMw/Sq2IoIIJ6sa++RRWAi9689z7t77jVTW1SQvTB8AnzRKo5ZxJ6k6BAex
ALnc80iiFlcYz6sOy+oIEDGl8bF557wLkdLbwDJH1t4e/Y3TUR0dgptYaRx2oUpo25TzuIJoAk3M
jZ7L/WjGpKd1/bgPuIua/tY0oNjoUBtpujQ4OZEsS4TW9Rn50cS8MRGNB3IDwPwLnRIqtuJDTqZq
EhXJkqAEjUnOvyTq5ejDNT7rTbx1BKm2l8QrObr803A2/F2fAcgfe/x891dQJJbfhPBmAep8QNLB
5vV3b02wkLzak0eDDUu6LEqrTkx8IvWZ7nrjzNseXz6OTBlG3UVN8weFG6UFI0UaGzQxYvWFo8yN
oP4hID9fWRvUablkdNXHjfig+nu21m1DRv3s5Kc78wGS+mjhN3YynmStg7m3g2dvkPFkwDnz5fEr
WgIMRmP0ihVwSnyOdFsBHjwl2ZJGNOnxJAyZoKeXwx3HWTZVXit7jJoVvUYWNgoicB2XWvi1Dfgx
Jn2KREgM0h5XAYchJK2Jnaj7VtDhSTH2kY5rHC0EU1cXBr7uatDRLiYtE1geFBYVfcX6xB5YzuH1
nrdOSA7faw2yNMe3TR4240RGTF1fLDXMn0GjwPdiGtzQe9gret3HuNkDEAeWhlEDf765nwZqW+Xa
+2nuMGtEo0hDd7CF5XEkTanP8ejBi8vYX5AuYl1hi295wSig8iD62fnOLqbX6/poT/gtOLnJGe9I
WAf/r2/FlPA6IpXRootoyUaQ4n92rKoQD9ZqIzVmq7zaJouoLdrilAfi81lDSAPPRD99t0lzpc7I
WWaG8Fv06GG9BNU/GpRjq4T73TwByc/sj7rPWNur41CPbRGviiXbjiw7XrB5ztdi+vVuGnvG9kAj
7xIDnd9Np4nEdVvlsgWYWD3iUe33rejNXXCKsQYQEYIMa3UkMLRKMS6jn2wwbqenrqyDcj/Gm2oz
94dbts2u+x5o49VAklB0u6dTCxZz4A2Bsr4yNW0z9TqeN/F3pK2EzfSNNl6pERrWGSkctMrUKWDf
O+zt4+UM70aRhfE19W7IzyNXwZe9tEA+ZMwDRk0kqQtR/dalFIRqj2CnSmIJD4clv45Z+l3y/aYy
5V6fhq7bdZMGlFt5BYMiGSMVK8/45VqGzF6kp7IVUizyEKDERqwOpzmMsOzYy5wVAvwS2JUlKEy+
9Z5gw7EwPyuQ3a0bLW2m92orofCv2SVitavv/UaZO0xH/hAwBa6A0WHGRXkdyuXP8tbFMBSV8dN3
KwO5AZ5Thi2X9EFUSfjLLXaJsO4kkW1b7N6iWVWuGJjMrZDKOLlgpth4bZeTvB5E2Pin6ynB7F0P
ObnPpJElE73EacqFXxhl6M1pZDkB7ciS8ZB3+jBiaHuylgmrPN89BIv2zayfjXD/IZ57pyJTqTQv
3tJ3wDUqKwKdJ4VumkizpnAs/hHkMJz988GMGpB1qXOvzNm6XNHuD9BlRqnqEiCFM/951STsEVH/
8XP4oeqpS72MIhoFtbppn4dMaZ1EhTPVj+xNh2UW+Lr7h4La1eWJC8MOgsTblqhmfTNHBMg9ANta
G6rUNUAXtALC563eQELADAJ4JjpXh4GznoCW97KsYnDMvNbM//EUIT38aFNCxPFibfjhvT6trtp6
1D9jwPSORAOzA93W65XUSB3RLmlzXWngylmx9aK99XaUcAoNBqNIwuOQpJqpD+rbWS8bGzI2le+H
J3/q2TTd0O4m7b1UkIqObvFBIdFxW9oFMvj2BXi6PjYtAp2pGdym5e92bEX7BRHiTjZGkW7+o+j0
1N3lPNp26y+LrfnsOjHaG1Tfsp4Up/5YnDGvliJjJrirYCZr0n1NPDL1DsssBbGo9VlENMSMm/es
bNcMfwvUPDmZBpQgjsztCikAitVSCQKFfzmMrK5cVfYtcr5J+wSxXlUpStoQg/8OlrEVVtOxjSN6
6Kljm3BwsR6788zmpiLLMqUBrsjJpl00fqXuK+Ko5+v6/uQ+V1Hvl901lyDR8G0kmCmDIVf+RUYf
wo7hbso2KCI5ivYaeKJn/QYNOe8huOEBhw1LxQ+FRUA9His8K6NKyfyHCE7acEb85EeP0yJD79sD
/gdvsPLSytTFrg2h3Emj4QXGkfWmN9dPBWUKYXalgkz5KF+B1SqB9inWtTASW1U2FZh7GJNmZlNc
1QqRvvPAMktwLwFUzviT4+rKT+ZwreLUxZ8Y9434KFM7cUoWI7f5sWC7aTTyIQRDcQZJ/YI1oK1m
swaW/OsoOJECY+dJowOLfdWfO6SOxyDS569FFpjVoVl9/7eiwjBajU0DeH2uxS5WP/NQKdw0UBZp
lix1GNBgwd1eh48jBjByU1hcOuj56Miyh+WSMZqzQIbTbmTm/rAoGgnbHDsVFubHLrsf4VJR4NIN
tPRbGWyumAhik0CJlshu9vFDdXnfA5iIfSaoBvffn3PgicrJgBiuugBCELJKh9Of8JRlJYReQRJW
nzq3eHNHOqSpefJwRmmlQKVtPppzsAsx2VEcdnRLruXgUsFv40PLUXKTku+8iF9PlnhALN1YnF0q
tsl3cWd2KyWCfZmnm/v4thvbML7mTWO7PeK8jcm5NT2/X50xVnLpXkA6Qkb32zSz8v/sB2wZCOja
GUVkFA/V2RXNEA0o3lMTE78ZYNAuwJdui8ljhoZ/Q6TNuKTj3GV20n1aSqCKPGSfPBJnIowNjKTu
hd2HFhHL7RQr6t0z5c72B4nNH6vSHCp8oSkOojC/kYkcYaZNjE7LgI7UjQLYksWIqrfUCQxUv0FV
ei5JX3J906SWeeNpEQ6gnxNvEEGsUz0nm00S+CKf3wcuaCfwfmYO6eyer/1k3+F84sNgbYI/Mq6f
7LeZC7vCwjxYrDnq/FKrLsluDmx3jbqFj/GavM85SaGKKtHk+DohPrdaL5m1xZVOhOalg/lee8iU
tV4/qvRbqvpaVHRNyYuzcy6adXS3KThjGl16vzH63ToMLXeCJAnGBQGn07wvPFeTATIY7kAnLjXk
A3Tx89uDGAA9D+AjzqLRqk6e96V74/1LyduUi4u/j8U3sZjK+03mQ2hAR5ClX5zzpDPeuN9sAHCe
vDqvsSBzE2miULcG10Rl3yL0Dir3XmSEhXY9S3bNWyiU/RA0eeDRSN1hQ1RqXQHPWLJilonscr/e
dTzmnBQRWx38w/4jtXhDig2oz+gKByuyqFqmiWMU4lj8at8bBqvCSuAOMt0hfh9YxFRS0KbQj8kQ
71rdw0t4rbJg9ZVzhe+CCsnnsDXtgk+GNTni4FENo3k2P4jMtLk9iyN+zmJuNchDtNAMggAnz38X
RV+E3C/K3xoVFcghvwQoCgi63A7kfpqLN8ituF5QZ1U7QR1Lid89WD+VN6yX6rKhvIzPNiIoKW6o
EiYN3+C03nM244fqudF1qBdU97DKCkDdrBS6WtAV28vU2VDVDT+YmoycX4RBi8HBDpVjkZhPsYcc
Y52Wo6j18ZH2tACxUyp/sj16oYVcaJR2ZTncvdnC12cu3HQ+oJT9jxwZL4EnPOM8W9atXIOH7AOC
7Z/HG9AK2Q2j8PJHVKPvTgPWF13Qk5eTfY8P8r0sNZ8pyk1mQHcqHIzPjvpnD/fxRonDSQblFoN2
QbmKhTaHp6fxXcFqDuHx8tfBn6ZVl17u76kdJZoByrSl4sNLkAy/sdNRFoY5qzsiKQlmR6kINrT5
rU17DVq+pZEQs7OvzETTrxXnSOoAz0JUrQNMm5K/BH/H1UdQkMVlFc9uWEvvS6/5oh+Qr1XhPnRP
lTPdgrL4wuaPnN0blkxOqm+TwJGM/4wxAV7P5Ij3fMAh7n1cXpMXvADC17DtJ9u7IDjcAFbtwHGI
pEChg0ZJk7jOtyAGRAMRNBDc9HJqmgoB6X+wVTilzanEWRK5ccXmtmhxcSdbJTeAL4Yc+Ybaxgdk
gKW7ZgVmTBPar+7dgh1zElyBFYpAukH04x6yUOTFZfyPn14Z0Z+pl31nj/CdK0QxTKIrubKQQnq2
iekFIyfcZEf1aNfdeSjlfUWAqVV/TlCFbd2uKXPuy/xMGrHfJ6+4KC9zQsptsc+BhOH2qOarjV5l
UTGAL8LA+ddtAb4c/Aq+4yi9LSuGln/z13OLMBSKSYPsUvWhp8TXOtp/W0vyRw+kIbEzuJS3VKPn
U0BcDrbLPYDm2cYLDE/srQa9CBYF5xAuw1dbU5+Pde2QJRe/Wef9JCMVmNH7rFZ/EW54UM+uFuhp
VUa50CwRJbWZ5JC1rGPAaszIGSgUfr8/niPwiBdzMiBejo+mjefjBN9uuN4aIA0591XYvF6v0nKi
c9kNvQ/ei++wAwWaHRDb3ttYHH03H9wXLsn0CCEUPDquylOQf00mV36zYRrkZpnPrOyaAHAVsD6r
vibfP71UEniszRQK47px8qldpXQ7zZ4s+FE7v07ZZPJSXFB0eOXtecFnC4DNXWl/2dnDFsR+oSOO
ksnkgh5B64yHFToo12MBCfCrZGWDfBrptVURh5sMHCDfQlrFFCF27UqJNRybHqb/qpAEOcYyzs6Y
Mh4IHELJGMXw+LF2B+49RuY6RUv2jHR8iqTJCW0GxZEI4L9DUf3KUL8/QcjoZpzbqgtHJojO6k0F
27tXhvRzPnb9jRZ6uv+8npHN5iP1B3daXUOpxxUav2PFStWNWi0GySAgObELm9jxJ05NFMbjgE+1
165YUZxnPlpRx/cesvNLY0MTIK+ecinBuJXCKNTGzMJd92FDtZAPuhqRhkwvnLeLyQedmdhxPtqN
jDBzsjg/VcQ/+IN56MXyELEj1HtrdZ5JTar1BFWqeUH7Wer7NVlpSE4pVWLqAqeIzUC6iNpWW/C7
17k57DCoFRK2TrDK14vmkAWVGUVGcLpHvUucMtiwqwk1fW8bWPC17cA7ukp0wVK9yOQr1djcnKEo
gwG2X8YnTvW7QooXit3xGPSZSdGk0meZq6WfqVRI+uEqwm6zE24o1sCKB6RSF6AR/p2sLrXGT2Pl
0Am3xgZp9c2M32lVMKO97+6REJ40Y2JLFQy1heHWrFQ6i7kMhAl801LSQdgbk+jHADneXXsGzOv0
QYgmu90srm2ITTKWuAlC7ZwyyqQonH2Ho8o9Rfvj3wUtx2uzxau8NwsxhgjdUoF3f6N+N2vHQEau
X6qd5auqy5LWYQrbLdHiB3IRzDpsiHY4NvciUJfFILLKgoDHeUoLjj+bWRgjlrtIfk3zBUqarQiL
YaK0w1LMqaffdR8cnW2oSlk8XLc75m+K4NuGu0Yc4KGIXeLE971KtAymOOzevHWX7y4ADB8hGpSZ
JEaFraN8wbPcDO1eiLJhMMPVkqh3nnmUwer8JSrm9AszgM2IZ+Kf3hjZVraQCrauShfuJVAM/GvN
U3CkZWz+A9HnjVriSKKjBsogSLlEKwEMsg+goVjjqghV9khOTpR6NsfpaIG1zuSuZ8VGtsZkeFy+
EDCfh2Wa/fAN/qsZY3fG/hhlpey9WPcL0Q559fow+G2/2SOyFlYk/Pf0ilXK/o2t9+0hEMQS0HZH
tXyzSKKWxi/fB1xtY5Uk8yyALHLsO5KVfZjVhm1dMQISp1/w2tjvtbohQLWtPEQM9139lIdT7WsG
hQK6kAO7nwh1AkkC7Sw0SVcp9vgRLUeKlFFKuUPOx7gSJUeb69n4kD0AxDUFrQU0d80A8kfptlf8
i22sl7mmdIHiEX5rvyz8zPQ0TnIGfv8lj5vbUKuiYXaovOOutDNVEpN//x5h4xwhGIaizuhLIc74
pVkBypoJ4gp/JXTJ+mVgcM0Z03I56mU9AxLS41LgKcVh/1qx1SGkGbghCQJSsaswwSI5sIAH7raA
zpxVJVDDKPhGn9pGFyAgo+dNTU6Pn0vcgKStyTJI/ZqhI2jydFgxevRxzrR1a080X30pp5eG6A7J
osCQpybxsYjrbJ4pFenOTsHWJ6HnB/K81dmxCcrzInduBSzWLHtnxG5Ql7rI1NaQ2/pwBbTv8cs6
8LKqz66qw8Vrri/XKtgwP4dWesjtj4MT9rrzIikjniwkM5sWYwRzwgEH+gI/OriYVdunGNzz9KZ0
i3agnSmh40npKUrE/jocuC3KWii4q4tQZCj7Q0FWle0hll0YiASLp0iyLBuBRPybKEIRNMUZKY/Q
s0iz0EyHUoJ1JttkIwZSnHPsySrUK0QbNasErii+2op96hgvlpylyTi7HAX0mAJOfZwDUixOMtYZ
gK75KXS2GWaDTPZtlZzx47ygxB11jNE50vb7zOqaFS4GvVO27s0y43Flr2JTiHQfIIcpWqQ34jp/
Aot3kQ29qwEUmtfq8wlkKs2EVn13S48gqxmJ0BHlhbOTrPoL8oWTA24Y4XAW/ccft78844+mBhEA
35Ql35pvw7ED702T+UqIvPGiYQFt54ahxdvxorLdugsr1o/6KCJ9yNn6JZCvMk/dcdHGVCKue19y
+37HvEmc3z2IJfBD+STyH/q6niGNSeYAIE4iBOCxG1jT+44U/7Fm2eIf09Spxrn1a8bWVTs0pmO0
4z4Ot7WzYynMbnboY25cdu/wTWO66qg3HOUuwYVh1USjHO9RtOifvpmKifyNdO4vwZfKcqGbq4p+
VXGnYp6qUCDQVkqR0Oh93nGhDCk3WZw0b7MlsINrurQjOgFXxCQBOwLXgIZr77AoLw6E7zk06G/c
p2RQzSYsqdWsmf+9bwRUksm6o2rzLXDZBC8wvhIoz3Zv3enUAj7IEXqmX6zF6A/9koRZE1gwM76H
uWReStfLl87ZET/5/K6KFaiX+fkSJN76CbCksrurzFcu9JN96X6Z8x3YFLXAiy8FbCzMLEAedYSm
aKluBLPPdepWXlf9Q4LVHB8zso/9sO6rE4ZnqZcDtpOU6YvXjctSa0Yr0d7Zky5XDMC3xGzCh29o
/F+ms5uQGwPt5RPeQsvABT2Dd+nKHft53lQ23KOzhWAZvsC3THLyyxSRIhW+QM3ZUCAB2fJCUXmC
+yRK+Cd9IjPmGxY74fsk7ALBqIeyYlpi8Vg1qeYeCg467JkTWMoY6Nl9pXEN1dxPMY5KtCbbm+Nu
mMc5IEixlC4uS9iT2OnRL+ScakM7yhL4j0D37lcM9N9DLlIii9oAJl1SHV3XTZhLYRqoj61UVoGv
O8wrkA3ORzlDE9HiYWp/4Vxuhzc4u6pMXvzEgxs5AogWuDEjc6IatArOfvvDENKQWnsD6hOWQHv1
ROgJPcujXRRvmc01vPdzOBNMASKhS2UZ4FYg2SvzOntx+p8uxCJciffayleIBESHM0qDvByY8q/N
KB+5E27bD9nUo7/FkQWDw5AxkGijWxyrO66KJhNCXaDU48BEuzfUUTdI2KtZWAdF7NX82GWicUQg
BlUWMLr2ZwUrLuEz5hKY0sOu2sNHbZV1vhsKXy4//vI3T9bcmVkHMyFSTA3KTruonrLYifwgoaHY
1qcVkpbnSsuefZcGcq0CQLCjGKOtTTjlB3PwCEkZfyMFrIyWVh0pQtmnKSs1qqkac2i5JyKFtxYO
Azlp7ABZDkes7Z71RJ6YyPQUCnOnNN6QYgZzLkTBaEqNr9AQ+tL6ERERLeBKDzhtAscLcAEAlAdl
HAMWo5HI7xs4XKkZ18vk8/ep6FNLad1bH0PjmP6Dd/AH+KiiAj/4cSrWdS53cyG+GWIhkwKlHNfp
qdkeM3/5TBYyT0KFrR5rI9K9d3Yap0G+LDtxyHN/8FKfbLpWXoJEBHrIOi06t9ZijcpWGTgJryFl
JJuhrsbozKvPvTbZoKs1KlHI/deUIeLNQ1a9GfpH65uGp/ZcUAdnU+2cbscNiZBWM3MfJB6stZo4
3jcoycvenFyUNlHRPhLCEwRbH6AfNYzvx1tZRc4PrncaqTEARsGEZHPeL5NLseHZwi5wdb9wtCGl
nHW36JkM9vlfEcosClA47MnaZK12O4Nfzud9qyy8bmtViE9fyJBWXzI51AgDuA14hlJuq4VXum/9
6Jzzi8383dMhYZ5TChUD5/5FGefUYzXNQH2TRNC2HJTtmmuUGYjugLq1L2Esdc3/WUKnyAodyebs
4NQ5/ug0Rk3bn9J1dbpxk/EZU4l5eSCXqVgs1Qi0kNnXAxDrrWbKQQmOPLZfXQgIBAj+JVg2Kj9e
hSFmSEVb4O+F+IxVKqhICdonY7E1uvCgf2og/L8K3hnxbHWInDYvK6QQ0s6Ub1X2izgitQ8fweSn
2iPl519L90qUudFzjddfU8LHzQ0G8C6Hn1TgqCaviUAEweCg2zxPzi3NrU1RNeIeHdO35FFNSVJw
JqP36KIu3fqA8HvpTksTtzFyN70VZDSbm0rchpSnf7CIEpo3O2DXW7mHg7t+Gt0XAHKnHEx3VrDu
PZvqZfQuqby7QJpSGR9ZF2FCdX7ABix9jarE+WjSj6eVyMkVQOF1PyNdvexdnJZSCr8/8M4IVd1w
DOenU1PJSJ7BUyrBA58J3kmRbR5GiWPoGadnk9wpFWWKxyAjkSLT/h9rLEbjgzfAIn87LyyQ4a7A
Acq8O07AoA+VqzziqN5xXDFkwW8XVYOOh9Tt8pLmw3ioDsLn2aBJBwaTzQ0NrdPmtoWwEtvl+3pU
XrNah5OGMVK7eHqfHMvvX8h4UMEauOtA0bQ3rDY711tSpr0QA8Nmj3fyN45YNnH160GSWE/VjO5F
S29it7sfUk5IlSjGptmHaLqAjQdvHMkQDc7GvxgpQDEgjIh9+lpLdOv3KDKUbVbJraRwTq0L3kZR
TwwGsqnEZPwP8AkY5HZDrFgl1WecXujuK87154vbhdHXqc4QaQWjGMzPNhu6hGiISi1Cy26URxoO
PzeSlgqC+OcOh5oz/YMfTTQSuK6lg4mL1EQDWrRtg0TMPNxZquJrHlErtyHYsqX9pS9ApOXCJeW/
pyZ5U58Hkafjy5eFp1hbTMdfWevQXY+tmIWz7lvZZEf4lNqYWPeN1tqTH2pNWvOONbXjpFKcrXRQ
8xN/LKeZ+IDNtoOFlHVuhITgPzC5E2qFTdn0YSSF4+LD/Bp0TRffvlZosBiFKKY4ULGo9p8AJCE7
7BjLMdMFBxXQvuCpyet+z6U/B59gXQgPqYmWRURc88m358TBIRb5M2slCnVR4pOQITJX4heVhISV
T9JitJP3yduxb8gm3i9QQzCCwM30mfcz1X6FSoQTyrTqEGbOV/Kc21gRpTfeajJ9qg6OHJjwWIqS
c04O3pYEFb5FfX5W6c81oq6eq6epdF+eyfP9E3SAtWfJaiqo/LyfC8UE+SSSiwIB9tysfu7j9k5l
seueO3wgiH54l/C1ILtD0sUf+ZC5GXGUzss4WycZm9Ia2GNlUHBq6xT4WojlCvE0ZQtrhxo98wIz
TOOJ8d97D6KQDzj4w1UJxIIBo1m6kFUGgzbWIq0OXhWihENJMXs634glGFaBlUnVyp91Kjsqe4cB
kNnnPuDlZf9uTNft5fDPuxYEk/9B+rT0JB/6ThCwXQQdTL4SvcGGtla8Uu01OdWuxTfSxxwl+cEv
FK4baXAd5A3C+QcJAwlHwp3+FgClhdhErSmxTR3U9mv1gEJVtCTTNlqMI4rLMz79JvCGKCFHyHEI
UPC/QrMD7Y+CLiqBUIE0hSsK4A3o2lFPGn2W5uYKbSkeU7yq6GA5D7zbV78DsVkL00O+L0sYhGT2
GWibACXS+o+z4zVuopParDlYLdp/OStebsrSte2cg3HETuZgMSAh3kNdQF7FlrYNetDHxcjbQzD0
UEyDW4ztIv8dsDe4KifBl9VgPL+z5iH8vBlOX9AWAG3ZXCE7KY5XL5h4twHhdj/dS9PGMA71bd7R
STuoyPRG/v/8WgxamLqHhOZ7IV8mfgXtuGaWjpa/Ni0B8Q8nCLfLAoZSfSgud4Q0HwBXSAbcLS14
rGFFVtBdSz3Dy+4hvSHcm2yba1tg+PcHREY9VMz/CLOX1AZjsvUd5Ifv9xBA70GY0sXBR2K90BH1
LEFaqlDV8hDkv47/TN5ap77goNsQptTP3eI03etypThH4JA9U4V6hSq+s8J125bHZBiC2f/8CVGb
7vsXGaV6tsFLipuo/e9JCDEZK2aRUbC+jChepJpwqsDSTqT4lrfgPrapospu4Y0wsCGR52I85EQv
X19UFPA7E1GEdVJQ2oC1YQKU3xV7MAtEmJ3jeDVaOcFuzVR5RZ0Rf5L9tvYzCg4Twb472KxYFrJp
RwUh0WjiZGVh1H523lJpmGyOh6SID637g3HpsVCLjZ5V/MlUcJ71WImZ+q9pTclakBuj+2ZhviMB
IkpHDIrlgKDw6GCPPciXOhVEm5kD4xkUAyRvnjwkuFWCpEmGrVgE7kFUzQA/Jy3yh6gMyrbiQByP
NecDZ7V93RNfR0q3CYulFcLrfkklbQ33+tSiQ3CzJpI2U/3YC3aP11SAeNlAQuBQko2fgRt+M5SC
9NSCOi5Wc3VN3LcF4U20mc0VePM9swfJdNqNwpQz10NNJ6G1oJ+wyUcUt6gSTxo8Q+QP0FztVzP9
YTl74IeOWFowXCkI3j2qxRJywP13SA865XtGyIxCwKDaJdvfQFAcgiawYfywRwOMaxuRUBYwWBo1
lz0hAJf/u8a2BZmjYo8rUNoTzcwFy43mKDUNvUjL9WIt9eGm8aAWykPlSISJwVeSMpt3I428B2mI
AgCVPPMIJsjDOecvuIku8aLxBUVEfk+cQmZho8OCX57XrVyl88JqhPmIf7DjgJRCL4/F7tR+McZA
dlgSap+Rjc/NGFFi+/RSOkg6h3ddIkz+UqzhHJ3ukEHMf1XBls8gJLPQiiwlPRooGCycp609nXZX
p51qTrWOfCO7ct/bGX2OK9A8wqJcFlHSz+QE2xihweBJLn3pJkB/3BKVgg0+tkLIwn05AZeYIef2
vRcD0kS69SLOcr0TVudF65ugd8DkgMYo3kCVxfaF6USWQD59/mHa2mcoZOqONRQBfa1v18R4KxtK
f/A0qZwyrXYKn+JJ6BKTy9jIQ2e4l3jAM1J72VJWiVuclKoA04v3fVLdmsAaHFbq9q2ZhSMBKfgB
sA+gJr3F/SYwek5B/YfsMuvHp3rx7s5DL1K6YddkX0rcWguERZrubRUMGSuRgoLP9xtVjip/a8Qg
2Bg/Qi+EaIDGiInKjsXeo7LKdZk0EjLlfiEF+UOhccO8aU6s5shkkunR+SBnWHcaRtiM2p7HV7aK
h9GfJG4X3lb5J7pdj0JFQsMNQ79f3kbcK2d/q8eqwY66K+2ZNtooynTpuIVn4tsCXgWxSouxKdNm
V+UQVZhAU/ilm6FxXNarpZk5ifglEBi1muaV3FGV8RkGdEjIjVyXi6pAOyyS1nX7ONeFgLYxH0BF
eee3m6+xAGO1D0Uw2JiRyEtIuKxd+MNiUdVjwDjByvX5h+qys0dW7DcyQ4jfD9OdTIgUfchsjNGx
86ZAGMbtWn8zC/Ts6G2YJUPVRH0JZT27RiY0uWqYuAUnWMb/DzRhG1JF4YQh+PFJy/CZ2khorrqf
7qq/tUaJ186bENbZHk8fo3QIJSj1KV2u3QAdZnoIrkQShqt/PTAH7frojtDJCoxI5QYKhtVwJMoP
6+ssmyZN9D6kJTOR8HSJk0STWhbm2yq8W2UOKOli9zvJHPPVD4J0fZOwkJWwZb7t3obNzHb8SElq
Zx+snDiGZDgv8d5aIpqEuNiTDX12AwOo1rQgp01hcEz4R1oK0zgFomrfyeSydBCb45liFBk1ivVI
S58CQXH34KymHHdLsorveYn1wQXlP9UeKb4UtXPnOqiSd2O4OEYk/QXfeEOuyeRVB4BAu2KWJ+t3
pBKXOfd2pbvxDOfNfACkyODnIAfbWcl13NyQCsIYZMGH1Mf/Nz/ySSoEX4N/3/B7pJyNhzhR+2ka
cGOpHDzwQObwiRqcWRaMoxGvz38HWLyaW/U+khjIJAjKoRjB6TpbmFumMzk9YQ7rviD8QkgNegWs
mZzw/WUrhx08k2eizzWKh3NQ7DqzOGbEIYkZqfTeSpjPDvDX+OFpxWts+J2Ss2uJCEsmhEYqWrYq
r9zgtGS6TND+g+SUJEW37f5ku06HgZIr5rXfEOdM/AtQ0SfAk+QYwKIrHGINIpFFo7ShsPV202ii
+Nr6paDS1y6pCXWmgJNOrF+IV4wa0XIDD8aRnwdugPBYC7+vZbeCP1HXK+z6M8el/r5a6FnP7OWu
LlhhBQ2bvrmmVpvsoPsihGhLQYi42Ei42BRkbv3WeQKXhXn8N7uD7wLo8MYWh1o12q9182C0zGKP
EAXkNvGzxNa9GId5BN0IJiQFvDt0GBG/3bfhcbpdqtDB4bIsLp7NS0/ImCwCsmVQfT5yjLe6F2p2
2Vbp3J9wUKVHMHpW7z0rfayvifhur5hdwKS/+XhImoBnIVqrk5DoTLvkYIVy2nt7GceX39HMJu7y
5XcC3Vr8We1Mu5xVxSbo1QWYQ1Nhg3ffD2UgWftUR2GsnQ1vSeRm2WBvpah/VqhipdJveA4uFYI0
yFdW6cjRLxkCEPvp7Gr+1b3k1Hgqc0ItaOZ3SEqdzXyI3+lpW9VvrdiOwqd8uuK897qwKnKsrEaL
ihL4krqJq/ljG6sg4SkCfqN6vYjP0v89p1PqgU4CYfELI0woizqoccXMDdSFqb1IKSX7zIMTYuHz
/NteqAUkHQ0IbFbCXWqywVA4hkmaShmfuM4DHrfCFQhTdyupPPXxJZ8O8aLlp9GnkqGrZTDfzbDk
51Q+o6PF8CAqnwv7cizpF448jUZYF7KpxmF68JPSeRps4OtvQhgIW3Bmugx+s98W6F0DNBrKUaLO
QmexslOYO5NM5ztGBY0FaHaAnayeYKI3NdNbMTfyHvvPvf++Tcf/OSyX1LllehijoxOH/Hj/YrPS
oT00vNvW4tVVEYa55PhR+cTTwXG4U2bjtBDXc95Jjcnb3xkePjJaestIdjOpqlPkJNRdrnAprqrh
YULREq9M+RGYyLmWdk2Fuia04VZ4upegZDLUSTxOaUu3CqnuCSvB81F24tGyWv46SCxEpR78hXV4
dR7LerM+QQQNApIEDB63WxmBTRBJ44eLMYWGhfVKjqx5EzYCpmdBPcPBJHQ76QCFnfIj9Qn/3KYR
L+9MlKpWf7vFKcm1UHCJ78SCctM1anr8VBV79mZ8wQhmpSkmjg71gZaO0jU96f3IZ8zjFhPtKgoP
eMDtSEQ/F/sbCuxg0lcUGHtM9tJ+vAY4HBYWqPc1miuZ/p7njmSLCiHjplaAm+Qj+caKdoOi1av7
QvSB+i7BRGvNU9cIXSIy0mMntxHZ0Xm+ZQR5dqv3ibtwORWf1ts1/EJTFREQi/IKTm3/X++t0f9p
toIAaIdP357ZjMGy1LmyYWIcN6y5sXe76Es4rJNUxkoZynqjVmDUYuhs6sFpL1jzKu1tY63G4zJ7
ALJuQtRVF+6sZhkkHezFWqBObi+1JoD6mwI8CHFy+UHuW2259UPIIBqjVAcbGLuIebIdtYbFG+yQ
ae8FIAZA4dxuQAUIQ/ZXhQVqrjRsS1BErX/hDIGlrcMtXr3AwbzTuLPtT6FDmMz0lSewbvyXOeqT
GLFaCVTYo+QMiohA0K014JvVaPs4FmWjO2oPCuMNX5VIiWhzpbzRbd65qygnZrNfaO+aCMF3Pqaq
psCopaZeN/iq2EL/X9H46IJYF1hTDVY8NOR2ICVdLGxsBdmsPFsMjv+MQ1Y1HPiq8aVujeTpI7s4
xiczdzXN31PLnnDa5eow4zGuI1iH7T1l2rurxqEhDt519g/B3mCeqLcxD/cjtc7xipFWItcZiSi1
J7pwQ3AcKrBZiNiwWqhGgUTD2kWXVPXorr9EamL3/BpRz8eJ7VQt5xiwh4ETqMgqL4EZkCCU+KIW
wbiuRaPWYbu10uHKJW6UL/77BtwVQZVv9eW6a/pnKk/yy/NeGufHRS1RSnU0ptEYSrGRo8+U6vlB
RgTtQWH2qpn454NOC7gjK3apHJStRrKXk1NwUPI0JOyORiGKnMREBHxW76FL2v15qHEVmYmZiUmP
CC40C5d2Hafl4DfYv7M6mTgOIia6SvbwW5yqXH5Yskn4rbXx5wRhOa1//jRdEDoFNm/UXGDEqlG/
2EBLSoYY5B9ODrcdKDkklRR/KrX8IG0+xyDFQapcPJ2qY9lES/BZoQgDqVOZQVn3ek0QN0ijySrB
HXo0OEk9n1aSCXLVyJo2EC4eotUch73nFambCmNfuPX2mV1dkUg4ngoxVQmYyT0QTcW7EUR1zBl1
rIAUgIeWA4H8VSqvScMh4tZkEXqPfqbF8vw77TmDQkp2OhU3IjsHVJ2F+c6myVy/1EL87PzQI/SL
AhinUgzTvZkXzGif4rQiui/mAqbLZkaz3EPVhlt6KxfR+EVXiMnuXWLGsEuIQeF0zkoUJPgeTtqn
iipT4nrqqx0tLvOCOldaOXsxWPoj7etAridBj0+gJoP5fdlDxvXI6qKBnWmMVduvEi93n51sC5as
NaLZmqwXsnGqEWir0hwoZUWXw0gHPyLT6f44LXs8sY6TMsJwqFO7mYrPgJ8NKsGGsfDOP1glTdWM
JTDJp+69jQljXPivjSavZX9M813PCpFtrwGqQaWlQa4VzU/0e7/VAuIe0xYoB6KkW3q6VuYutBOm
DBCvdoJpC19OARJBc6/Lzo3Wk0bN03q4R8i2dg9QX/Lhy1Lmi4GCmXaLSB1tMAYsjHrg75BtkVlI
/sU51IW3TZWfirWe+q5W+dEVws0jyq3gVG1Qg+/7isU=
`pragma protect end_protected
