// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1.1
// ALTERA_TIMESTAMP:Tue Jan 20 08:33:54 PST 2015
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b2ekUi362riomQCdoRukBvXQYerJgAat+NOe2CPjyM4v08kCGJemfiUyrn+MpVcZ
2DmZO7Wwb8WQ9VBrqX2JT9tGkrYmByl/O4CIsp0x/NKrVixIRgqXrcg6wai4yg9N
SEzAyFlOO5nRwiFFw69Td+tc+vAR8SJwVI4H1uFmy7Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21328)
cZFxhbF/x2x0/KAy0I42BEjfr+7CS1vUcT1S6jL4KSAR9JZ5E+OfuASkX6bLp1wm
GTfDYLbskydsjSlZYGWoc9hu5iVUOpYC0YBLeODnwQyde2ZQXoR9ApU9pCIo4qHV
MJf4W6tFWEV49Der5jaBqJiFgi6QSi8Kna+Sle/XRa2QA2GU5eV59dDo5szHoskp
HaQY8E6MkC3chV0C9dj1wFMfa17CzAH39iiDL6o2vVEUpC4nIenw0027e3qjSXwq
VakY0tWMKVSP/BlvtkX3YAbm+An3NLEU3cTnfV77V5wlxY4d/VwNFZ9WfbF3paW0
fX4y9SbPQnF3xb67zhXz+bp4l8t2GdMmd+oHrqub1+nf/B5SLEqjKexJCc4K+lw2
s5oY0iD1UxubB8e0ZwLT0atN2LpeO47DXZ9NPhEu5fjfSzg3QKw6K4vAcIE2DOAa
hhRyEscbktUKistdtnLbUO07Czs4JMWQ1qQJZS35oucFTn3lfre/fNlMuG4SW67z
rzGJ+8M1qZ2uEvUbs4FBKjl0GPcwu8hWJgoswIp2NFwIRWiBd91rjmw1IgcNyroL
/Zc50C9xZBKQJnYbOYaf9xst3pjnw2USToLwcSJTUPyJcD5h/2vRoBnpwKuNMVFG
NcGRlmsHnOUrwyBgr8Fd2PZdhQe/tTKNETxq9iB+hAyhTDMDdLTyBjapwb2jqNWl
zrtVGpF1O+2QwOnhC8lIu2yEMSMhMHLxLdNjJniWoQUeDYUlY8IWRqWDxRcX79ok
JvE4q97Oz0ayUAp/zFFzun2mmnvWp9A3QPuGapsfSOiXl+l3mlYAecB6wG736IIJ
AUf7s3OfdINiwtZvVLWaUa04KvBFebGDZFEjP2VwAq3zsuVkzqme4rc957Fxl8RP
Xd/ZB/fQrFnEsm+MwEnF5sad7MN85nkHOec4HFoxzwsuHEqhQuUIUJmpYHskcOuJ
cGKgddj1Q8BS7jJEXRVAqjNDm+0u9jWpVMcbMsw0OUr2iq9jS5s8vmyfl4SvGbN2
7XpsQtWxLHQa2HcCsJ57dJy2ZgzEufBLx/kG24cfUc0QtCM6UOVwhZhDrAhQ5Iwf
vJynxGlV+87g5ViMuAe0E0uLQrCgwVDQlLeE/ZiCqPrHXvq/JnA06TnDlboIzStZ
6a7hV4L8HHtpjQw3DWmjV4E2Sbltj5aH0c8Qj5SKxTBVoPMEMxXCHKVmOnf1ZwRY
2nlznRXHtGxRr9QvB3xlXWBn/S0ppBYqlC3dNEIgy+yhs/EZzG3gE3qJ8Z6LQDP3
CgyYIbXPH34luAWsDpch+4ujKKJrbcwhqrCK4Xy61+yBGaeKevCfhNL/ggoVziZu
JSMA3rurxCTl0iAfOSw2aHQ/EnCrK9BkpvaxxWxCm/lISBKfsiAsu5sSYCFE/mQJ
atEcVX6SbSj3zAkqTuVKjrHe5kSS3SzpbezJbxVAPhpyq1TE454pm51LR/Zl7HBW
vFTWsbDcWhCxSf7Z66cFJYFsUJ3ob5wtyqS93hORO7KheVNTJmXVNbY/+mh2gm6f
gnWonhmGwRgGUJYADgqFLKiyNGc/Fwj5uZbzhgodLOKElYw1PucvC11BjbUcS7Pt
wGCmHYVn+KWzPH3klPh535h9GkGP7NVeHX5woeNQ1y5y7pp7A07NsqKobLd8ZG53
msBV/Zh1G9FWfn7zJRCgyLNI5Bnb5egmB0gx7Es3AopRmK9+q5zoGfQ0fOHkatEn
krg30WHzUn/VnmhCCBxzC1N0aKPHJGLwqRdtG+dzwAj9kzIsKyrzLfsqHizXvQ5L
oWoiu/M8j9yIdiUsKMLVpbPPw6QgLW1/DABrZK5wcYAt/OjqYu1Pj2hBO+wFnbEc
7NsbqS9B9GrpB3xjh2ULneyIjZ4iNABgiPIZ6WCJgO9+xscXt/LoBb8gBYe+KYCR
TpOdst+91tVCys4Ve4t4IluU65UkK0PBJeIuO99JMO7ra2MIUbIpaHfuFR58fr8s
dAYHrLo0usuYwBqKAUJZ95NPtth8LY2hvlLebi/h0bH98jqK7X0tZzzmpu4SgC7n
D08un2VUNURgOAHVbXMyyDY0+FennDNMeIOUqCrh16RnVhXtvzzkPMmeP9/szxEm
8rMOhrF6AiI1LkOmG0xB7KJ8vXn9iRSPV8pAy7Ks4S04Cjf+fajaomDYOzDAMFjK
wqqomn7ig8X22WtjF7aeduD7bluZT/64fAqbNXPKooZDpLDl3JSp5pJl2I+yqbyN
rs/ijvI+QbZyj8Ny1RBGoQkIUlgCd4pWYjKW+hbT+yicPMfnkq97L5HlB2OAH9gV
UI2lyeWKI19t97I/jG0wcFX+qI7OjqLi5JPl8CqYaz6rjELnw4G1X2O/SOoxSogm
/RISFVzsG/kQ//EdzgDyea9URHvrpUK1aplTSYHhsIHyNi7RRcZKV8wCTakAyZEj
GoYP0mHh7T597Z08q9uOJscmKWb6cw042JthMn5bCuZHv96Ax6gcQkAouAXPwrY3
knfdAb7wCZNjWLBYCDL1P7fcg5G6kDcIDXAOb2sAKIq1bkEalDj3093BOqGDj1oW
GYVMZbpd5ZODijLCd+Op1+B4h4hphoplaI/fOMDZQCD4IwMXJ/hD2vC29pvgcF3X
ytiSyLn+6p/8rlWOYVjZgvbKrR0okGMpTzTuF9kZDxyDZEKLML11g7eINpBna8T9
/c95Q4WTJsrAFHKYtRxhnVQmiCrFZFwG4oZ/cgDM6mu8EmJDSJtvn0vz/WMgwMa5
H4zqwUGw5UDXdOzNSKo3PTULcYwVuhOJF6qyhiQwVI5T4PqBiTfb5L2Ck/wBaJPU
2e3JHQ5G3Thp11epimI886Tx9ne9d3lqvBt9jo4HYWiv+KI6r0k/C7UTH6xfQ1Z6
81eW8gz9d35OKxs1mJqjO6xX4lh/4a9bQStKT4UT3sYTMl+BFlmrtyfiBUq2pL08
zukJqbJb35I8JAGYy4W68iUPbrml29c48ubspDG9+NmD3xYzOD3a9lwgmHA0ccVE
2yLU494uWspnhCgGtPK25utFeNKqeJs1D0ZJOR89umVXknHpUweSNsFHulvBgAcA
aNZd34RhJX1eJYWpYVL/mHRZdD8JzTWZNBuyvoIi+gKfkcI5pSD5hCn6e840kMwR
GOkYUWqX604CVOd9xdVL/RevoJrhebz0aZahq68dwBMRhesTcC2/VbQp/gAXhCa0
aWCFYfAJCR+N/NULL4m1rhDk9eDwfs5/yrx2EPaGSLHo9vrazJfzpgOHDwnF8haO
e61GbNh3PZpZNX4WLD7g2ZK5mVQFTGRDhWOY6GwVuNagvdxHg9Agz5M1TCA6Uy+N
QRU5kvSJJ/SogJOwB9bx3c+hTB/oWgqHUylHXEPBYGwkv8VOyjRmBPJjY/Kq6gew
WXZiMiovUTaoqLc2q3OwGxMT1RyI238vWGJhdYI1HivDHrdxsofcQlluamTDe1j/
ZA4KMWsA/2amOqnALxWpwElWbiXDfSbk7SOL1dVa8PGvvrW7ndeC043VycdEUtIw
Fg8Ffp/jSHHREGOcN+b0q/PmvPY6PuJg4fADe+SJmUqoqooJE/urj89GFFlBW8wd
xL5WZL3jzxMSwEM17YL3sSUvngGUGyUhDuRDIjFOpDBYyc/VOpJtCOYxaspMqG07
G4W90xBsSL9DIwczkPFs/5o9YUbVR4LiTySDKpP0u6k+w2xLJcEEjOy3BFI1VYOE
OSY0rF/SknAvsyQgYFAL3lxGXfDReRPrfQ+hhvCsk+YW4UCQo6fbN3g4NyaAzT8P
H9JRbspuv1jti8MssR6J+vCTbceYdltdB255k79Rr2uUIRjpmHi5tMV+wFaHIBId
4cUpRbFbAOza9P/SpBOle5qmUwiq6dc0dkIrrEes4cI1OKNrlshPibk43EEzileR
Rp8bMpgmFVTb1yHz3msBQhyIFQfNI0eSz5MCZfKIw4x3mkHhErGJ2F6pEjm4NqRV
C+80tLFzTNhuhzqoQqHsRmy2mhM4vFLXnr6e8iTsDFOz8gPOzmlu+VAymQG8PBnm
R5UmrHhhJSjIFBHtkObP659ie4vM1LOxNPngity5aA1RIELBdEmLXg6ILJAX1dcF
r4hEMIbMvgZaxsK51xruIlJIX6LASFUKD7GTO/OgkXbQPDVxxHGiZ4e+VezctjyK
O6l6dpxdcB7fgobuB9zTyIAta2QZZUEGYdgZl3VDYPqH0VxhDCAmJynlLIfx2oK2
456r5qVzzx80rysely8fdIDI9AYk8aFfXJhDQ/Z3P+kAYiGQRt9qrtbQuKd8Vy6Z
OGcFfNUA72i4oRgizdmMm2mwDoEhzcq6w6DQSXx8QSnKaEjvsWPs2A7jtSqelpDR
Ia6uhLn03QNvOfeFX4tlZ/EcEoQc3rsNkWLcENVJ+W3bDQGi2xO5J8FjCiW5V2o3
3wxFYE14bAukWGAkcNwmcHbDINQA+1n3QUFRhBQdsSsAOcEx4sXjJx3MO4LNz4Y/
9O3LpmtSJwNZ6qmu8YQ74zDLWHTJHp+KtzmF/KbxxrksG8sCHB62QCwO4Yv4duZe
psDgSA1+N4kFwSX0923810m3YXsQhOR22XHQ3UwlnnFzAz5dVos2BpyuuZRxAAOx
BqHnDoTKJ2kN8BSvO3G5LXUug+4RNkBhbb50Cv+HGRGkb5GYDraYbjj7n3C0DsNP
uDMJcnnF3TBSI4+OurG6pSappmrr5l4gBA+kATuQ+UGfuaRDvMA+E2CQqj8JkCRI
TIMYa694CIrkcbX8R3HKpFcbDgt7fHqqvQOudp4GAAAl+Ne3yEa1sHl1YEyqANhW
vnXlo9BBgeggEUPGrTaG83BnpXccauwjL1FrTvzKHjohcg1kpdWuoi6ZttLGd8Nt
g3YAZo1txq0vUh0wiQPPiih136xA/obp8wGCI0G2QkthdL1vqDNCf7OU63iPAyjV
JH9wSLNm9W8jIvXR1qfeoXuGaIj4PsWiFY/TULTjoUP9ZeOfbCEBJY/4oR7GKHUn
0it4Ddh0ET+XlOCaiTUraX+S/ctUpKXDd90H/nVmT1AqfhQL6Y6AwVNqojU/CEV/
TtpkHc0iXqBbCpx5qJai2mpeEH7OK6/PYkSWmYQEG66wYhlqcRlBEjq8VmGABwmU
tVijZarbsv7B7AqyZgnHrSEqgLyvNhWrPBdLOK6PFWH0pY3enaNRtTUgNrBaj2i9
efETbCftkmR5mlKYcMvVLyDJ3KcF9Jqm7ttOIoB1f/e6kGWq/jqHh0Aupsk5nlK1
6EKdGm5kTyMo02jrKjm7afpfwThCEQztk5UgjIfdHrZ/h9p5i2FX+MYZmXVyIShu
qWCnJnLUGkXLTCcLzGvaBzJVz5Lb/7HF1wz1dctKIQPm5Yv/Egha1+X+N574DVg4
NGAqG/c7X7CVH8bhan8hfxIzXslOe5Adw58263gsjjO62E3yG1dtg0xe/+xqhVrW
DVSv0eqJiECQP88k+zJ9MHR2vNAhqFsLwjijHgTc0o5se+eoPT6r+5wNE1UF5YpK
PI9grDEqrTCkJToD741X/x0YkX29BQOF90tshhX8jTwx2C10fKbM1CfdyPZa7oco
qtJm2hQUQwUFInRTBxE8rBbCQ8MSXIP+0PBWK8pdD19ITvfSVR0MqXYy2i72ZGXr
hVl5MNXb0B/92hglmSf3liRXLjXiAkyn17xw3m6BYkgtXXOQy8HDXmKvDS9CDNS9
HNSgX32hZtzQl3ihDBMUwElKra2dw5PCIORM2df1m7fenYV5IY8Ozlf67Y1/gU1W
VgubYCbdBm796Bm0uyTw2d0uEpYi5CZcAWHg9+DoNGAWzVsT7RCmuus/mbNyGWme
/OTUZuZFSqEBYMIB6bo6/0fi05Kj6BKX0hC0l309TsWCXxh+1A6xkL1F8zI66X4C
aJUaYb53ype3xI+hcVnDSEvioqcDWpkbcsdLmVhgYa0AAppDFSlpCbbebbmddROJ
81tYpa31jwbP18oarFit6GpMITRlo4eoROp9TkZIVBZzrYsBJfnv/0BCyjXr1Hft
Ib+SdJ/2PFrDIibB6pO4WE1URMii0D25MDRu9LV9NSpmqGj/X2jAtGU7YRTmFNtd
+7KVd3/xsnkgl14cMejUneFbmF3ucXeI3eO+k7nlmoe1zvMaOMOT9ox7+QZfQ2nK
RzGAEfzw2ltzcB0h4H/gSdB4UZJaUq5DJwWy85OITjn3wahhe7b0LpFyLSuSyjkM
bk9t2YVpY7rxDUWi7jlFnvaKZ9hDv6FSMu+5ykuDO0dOKUDaKfhYLo+TooBCurah
5hJrQW+D3j8R2N1Z4VRO7MvjQWm/QqHmsgoutHD2CnRX+hGB9Q+IWWDgSfU9sge5
l/RmxPU5SZFcRxn0N+i/ib2s/LlcQMzFkkZjRymYp6gPywEI5yXdAghbFga7Wrkc
60FCzN3jD0imCjbxhGVVuXtjQjhUtXIguYaSuYs/WvoBJuI3QUBpL6iVY4RHYNZV
vTtBEhO7ptK+onPnFbmL7P9c/KMew+m+BBwDt2F1fz+PEH/ZYjw104bbck+SHxCI
Ayy//xRNUkG6TPfrWknU+x8Xx5u6NBNBUOaGQaVn/9fPJ3gwVbysoiwdmrvzhDDN
tUYWfbnKRAHA1WMNuS16ZfJ8us9DG931Qs0BNAqPAdG8qbe6BXhWzxhReHSF0DmC
T4u5sUkLsIs/DKlvwolZIsIrwhmA/oxD1NI3YSAo0HQHFx/HyRyFzcRkrRxTOsLC
zO3uvo2MvBZqQ5/MZHG1jl3BOxZsep+g0lj0NPK/aYec2eWZAaXzUY/KrOsDAlsn
SegOQW/fhUzUsrLdZsIP4Mbfv9i6pHpDAwEXN200l/9FE4/juBzFEOfrfxMe4YAL
oGubN97yg9gE6vJbnBV2qe2nZO88Xqe7aK8lUw9DkahSnlRa/ipWVEle8DNr6Y62
f1IYAvNDjRaLx/iUSEhbgn0/9Tx880o1XsG0AHa1af6Pc+9KW7hLAwbIyH0dPTdA
YF1l/bb9ofwOi39k0AIa5aEY4KYizG6uVLrKn37Ntx7Xfd36jhMmKPYiUavDi6Fx
zA0ITQkByIKNqQTBNc83lmi1v+Wj3FSzAsvnDWB726nZKZQ16nvZe/RW/CCC/B4P
meJFsz/APDehYFaFrsC+rz6QiiEFeWG/pScA2VZ3C1qpsnH36w0rBR97Grq6nTre
XYvMjkGYT0AVIuSXW4U56N425P+o+hIIjK1Y8j4xYDn4jkmJZSZjZQ1IMrDbHdzj
xBKl54GbuILKTqlRvPdzdgde81dfXOQ5uEXNQqj6Zb6mAikOd0UiEFzJNWwiBB1l
DyCvhHTP/Q+a9ueSYXzetK/JPqMYD1xNx6J2yEvkCLsehrzftBcQ0Yw2VOmr9u2K
LACycdndMaRXu3uK684/lFWW8CxZZb17+bYaUobnWi2/BYbs5O7c27blL+GS6ZRe
mfAY6RzZwtlRinHPo/zzcXmV0+0sz5q1xwLIdd0mtLs9/E54dt/cevL9uJRW7x0s
zatr5/ZefEfGZIY4MLlXERXZAl4woY3qnvOGekMHg8A0bPfBHkv9tM95FOQBvjcB
ktx/JPCtzo8+6DPgcFErwJyw6ivzfaNSSOMGSL4OWIqKXALEI/cI8EChKIKhcb6A
UjVT5f3K6FuNUSOuEdwNnBmRdDDwidzzI5y8RKJS+/E6bg6R4dcvsQaceCKPCKSg
vTecf+NLCuQ9gikxvN+FU2qSyuG7m+dyI9Ai7AwRa3FmdLUuTIvZSve0xDb8LbCu
vUSxXXcSfIVaxDaYhIR+VSDu4f+e/OOG/U6o+5TLf0flG0wAgyEH8xGIiZYvw7gU
+KzwOhbRXgxrozG7q8i7SueUz0VeOqd1+q5wDXOSpcgIYt6eegEQLXeYE6P/d1ry
yC+0NnVn1v472xMReON51zMpkO3U8Qx0iYUOqpx1iI4xpe2A9CqsA42d+S5E1TlK
mT3STmmd1vWO/oBXCFz47Ilw43kJact01AIr5Kgce/9phWOQ+vmZxIkbDe2lg331
b5ca6sPNf/LTbJ17+hsACca9cY8vOWTpjNWNNE2QpComNgK1eB7Y+7gAulyX3qLw
KA+ordrsFSx6uNhChew+O3DO1lFZF86TVHYwHuknTj7aY14Z/8TZNNcZuA8glq1l
sCktZmpx/Y9cfvgBldU8q0QrWV5dFbQGGsNA8rrUi7JPKEguqLLsw1vz3lhUbSdd
HfmyhPvIEbAeagPZA0cKeIPcylNXA4neNxmd/6LdJTmqKH9KMyf1uSEd4haakEU+
WiBQ3R/k+QsTGi5jaQH9RULfxOUSZUJ/dX7hSQShT+hVt6WgIK+Ohepo9+yPIVhS
8Znx2E9fTxAnwKZ3Ty9vex5Hd9B5iyOBuqB+/gMX+2kQah8BJouiuXa3rF7tvX4C
UXYlXq/8h78YDZZIQiUlFR1XJCAkekwoWU5GEWsEkHjSvGVxnT2RWOh0OK82s7b3
OaXYYRbgj1dt/7AkmtDni1vYAvgrDINeko9TNHJRWicul0kZCzUnYtSFz8GMhTow
dG2/6NjxaSC45fgkLnCzpz+Zf9gyAcyGJ5U5oVqycHRKLD+ffql4YosCuOGiNwEe
aQr3J1J17KWo2X3YDATWNpqJwiMuM3DxWo7JnewHGPSum6OWkHEy5Vfeq0WjGwLj
/2s0c++NwPRm20GrDHkjQlqUyjJhtQY2Sf5L5O1gJeI59HcPmX1MI1OHRB3FMNse
yP/BnYr5Shja2MgcIgAkw+4M6U//26gva0R3rODu3O0S9JQj7Cht1Fkuq1AydZky
04p5vqZxQtSvSzae0zHFIAYsxf2IdRMnRyKx0+sogISSHd3/r7w0n4ymyyg/lSE8
59kTYztRb4BvwqeC39aM3UmSpdb/2BqM9OXgXLKeUGYfJI1umkXVvi+rOc2NJjb9
arH+uUVvVamPYmJoa65h6fiiXrb965PuNjHr73D4P47VtHiz8Aq360LovEzeVnOt
/AYnbviMeCGNYBnf+g+KcqMMQ8+vePamDccLpydrGfMo74PmPlika902W7KmOwpj
Jco64BPjihoQoUxFAhZj0U80K1Ud3orFKuxZm4FHG/cxQGqGVN93wpiBsvEEn3+w
BLsesAeRDrF8xe7tYn/r2RpnjAmB/pVsdZzQJXs2IkvbVTy2qKnSkWDwoFq1xm81
R+6j1SRTnTfzK3rJm+c87FzAZmygWbkAjIATErfStVj8p31O0GTDE2jRbvRvOT7e
ATulcI+kBhjeLFd25LTalXvIrAWY6iAaNjEFsrZfTPFSDwGKcGBuf17sPVlsDbs4
9WZJelBtBabuY4JzezpNimGF/6UnL9C5PxgIyF438Vmye67yCB6QgH6ntm1nJBMu
ZoSNf7UWZXqf2cUFhL+pPLXlWH+bbahkBdWNVhcJP89bR9XaOUHedmZujDmbgIIW
WKzRY/qXeNqpTE7HksfzLSoXMHZD0FfP90APgKhyFKf6r8NxopHGbuNWyU/5UjaC
IAUP/4pS7u9HqK+UHND1yK2ATeYaVFlZfwuUkLeGVFF3J7EshkcOrj+AqCiSOlwp
FN5AekdTYPFPc8wWJrNwGfo13d6csaKdly7bHHoLXL9MN2k1L3sEMaVxKXh1F/+X
Hrz9l+RWAI0/HFR2zwMOJ7rG8eoYTZHXCLT1tqx4dWQOhkrtrYLLbKFPXgSa5qrg
pfdj0dptGP+ySjzG5VwUj1oNBCw4VC/3Ow83KxLfN1P49HUm8JMJFOPv2wq06mxF
8RjYS5sN8UxLWam1/GmYLRK1Ni9e0IGSOl8vB2XAysTfwUJmT3F8sAiNiBjjwRM7
d4KgXJqyjiNGH/XT+fDhX/k8aAvk8SRreD3ErkFp3Oh05bA8JdMopmFBkMJHFTBI
0JARx4n1Dz56O+IXLh3456242J/RMQBFaDvlhxdiKkwZRaWz82URmHt6k9Fvv968
TsVy2VUtOOg+q1cjUBcKJ5rHr3T56LM61kNdJisfhSbR1tzi6P3OCgKCBuwvIH0I
noVf68XWF7yhw+/dpC87n3nJrGCuzMCSDHg/8maxdIbbeeZQHvdG1ytCWXjaovfo
738CfAZrfJhVmlf1SEKyEpta3QyVm3Bc31CvdMq0gda0vFMLehT/Zsha6u+ODPBP
gwGEYY8gSqUprCIsah6rCU7wTpkhfiHGSKeOXjsja0CzBXNVqr/72gr95/0tEqIS
tUWADv807RuTSLuZ4KzKxilrZj+r/gcnj/dOCbIrRrwqdViW0HrEcLRyHq3pinT3
QDwef//XhLkqNnRMKPRHvlZvOpLpqxLXdvHkoE2nrKEDBMyjrg2ukKF2HKnZckHj
fPHOoyAPl1E0tSXNE2ZaZeRMQjA1G0qLm/GM+L9TFR+wrY8Z7eQPfh0jHcNmsfHp
bPYduZB4mNDhCMrm2kNeRf/Ulq2uxL8z9EPua4R4GzZDNxp1CDDzKV+QjmhYrpOQ
YdeIsgPVO9l5FZoX8GTWmpnLrQLtqGdWTSTxFjSzzhIw2jEw6I7mLtqv4oRdhVdg
BHQDwhCteKcQgGX0bu/crPAJfEzkLcIFoZRcqrmrBppu/XEti63tKPtVSlB4P5RQ
uLEOPbhLgTZMXvGLkSf7r/R6X9NNrs5vz8RroZ4xXGk4IAGcVk7CD+t4FCiDa18F
ZxXEYTWlZDkmNqH6Ire0KzgId+NyCxlkM9LFxRYRHhCJnlQnjMzF74blsjhR1cFi
lo8UKnjBVGTe/+V5rCn7EKf+c6JukpASTcPWqdrdi0utVygECmBW1aqH8WogIhB2
KKyIXlbC6mdpqmlytFNC+OKHOkgiAK3b/k14xUxX1jkK5Dyy/d9m4kO+AzOtlCYU
ayt4KnQiOPigYGKKI9alYdqE7/4jBoHVZ6eT1C/RdTUK+T9+OK2fNdQTjG8xd9EV
MJ2FSWVrtx/Od+0N9C1kqidHU4DrZ02N64nWVZ+B+KseSTVdh2SEwQXn6pgFMseo
e+IpH0WBmIG6XgfJZLTCr56+gzlkvdHyjc0hltNoX540gVzwEtrbD39PZFYkOFT8
QdRPNigSwJXkrSnbbmJ1WOmc/OysspRpyxoDNG0BSaop0PjaACt/W6GITwPzVJAT
RXK/ZcZjTcbK2+XUygu4tUoH++Hr6jk/AXfAE0f5AGJCcn8+9syJ53Eow/NxsIXJ
/E6UYdQHh+VSvFPaSlRVmDoUB36webx+p+BUACSn3VmxYRMWGribcY0dkUgOwRMU
HrDbZy6Bm16luX8bDi/UAtzA5YbWZvjj+vkrquLDhKXe7GzBAO3clpDCzowIxCLY
5hShu7JEX8HNL1EN1tqviRcNuXtR8pSL6C2T++JX+yPVzTT3fVuFHMsznSRZGAxh
l6YWN64/DKC7Dhy/nzPSfzMq5vC/3c4CqImfNEKaYLON41tgUFo0R7aYhAnA2jQS
5HP/L06FXC6kUD5TAs/vtURG6nCwi0aUYgPyIefdTMxeKOltljhAr1iAepwLBRue
SjA/QlfHzx5Fpr6QnNDMTYpXBU64jSV4CfztLSPZaN9L4bXSUBYi+aefQKjFL4On
vF1Qn0xe+iO5eCs3jc5HEPMIgNa5UdN/mG9jaak9Yq2t4qvcg7xjZ4+ib1ALBHJM
IddS4okIaUj3P7Rw2054b5yD2tbYPKI3zSwWfqH5IacTXLXPcUkvCRyB+S3K3E5p
dSn8j0l8cD4nF50LK/n/SeF2qodtYtx7f1cNGd9XMgXk76eipnfXBMO9WIdVoZAT
9NcbyC1MCh4IA6Q+7/180eDemw4wMAmpKya8gQTN8BByf5cDp01MxhIbeN1VAIWU
5wslPKJn+Lt6VSeXCyjbSUMGWWjS6aH/0iA43qgXeOb9pK6mLEt6MTgNIOYqUgNI
Jxwy38bGss94tRKFGEDKuqc9gtVHd5dlfY40tlLW5eeFujf3CSvJ606sww74tJhG
WGAmqDWfIsRaeVq38Y4slUJaYiA3J7BhXNwdusItuYpNUzKfH/pqdlGzw4rKSZ0d
IHjnNW3b48BfWl2TDsdgljZmxTvhp0zO1BXpHVa41NS7VnihsxObh+O/4cQzll6C
8xTDBtvrLIywpctcN9Yh90RhvzmYhXY4t3qoKcAa4LxQUt5xzDMlj/Suh0sv8E13
HkvaRV7nTCVjb7r1+GOTj2zX04suS054Vboqk9Tdf5EZpVN07h9CsJ8J5ZneiJcK
6lzW6WXrkrne4jslWK5ZdWpfZ+d6pnNER001RC7owXV6JVaPobBQ4nUXubBoa5T0
IixHNXKYECBn6WiRfNDQclPhzKIYzI/PrBldHml5JBioNPNzPkzMA8zpNA3lUkEq
r4FCPHfXYmg2YDpyuRREgFMJBBPpba+QID0OrDPR7R7JdnP9f7qfI//E5rXVnd2H
B8gM8jHyAw6qAcKqahTcB3xapHkbFaNyNYGOV7cJnkckAcUrT+r0LNhgdLsPrF1b
DyzeVVRd3lOuyNITt8FZFF/wgQZ2htcszxnI2HLMVEni2ce6dKb7t6grhMeaJMT6
7jskm1eesb1nnbr+czAjP9pYWcnVcon4Q6WwSjfdDd90hO7TZa07c0BHKd9VMC66
bN5/bzMCLYm7hi1PCPwtgQXgxOpR7a1CbXBplAMujfg7zXwsFwDJMrRkbuMq7V7t
nCasvixlfXxt7GIeRbMYySIGDa7/Gz8oy6Mg4Ue6AgVcx3wCoDSTAQ3TgYMwBtAr
afWQpSP22cdRjdYG7N3b/YoPgZxyym3IzeS7stWoyODO0lBYbaw36FDqiIhZ9YYx
bBVfTPUNk+37bW4DINBH8Kn63Grik6ArxTvB2AT0UUJWDHVZ+AQ5KNAI+HC+uoeJ
maMFu/WPtBXv8U3hn5mTPt33bAw5dWtAh5LXvurjJpibMj0ROe8aTxbpAybN5n/m
V111DuDCPVC3Hkb0GUo9r8/7chK+MBdRC1lwpUckl4NSSB1TkSyuUyXf1XklM0z/
/q68l5a4XELFsUzbJsYGy1I8x4CB5/bRkXsozO4irdH7M7KyQgPcl+XLXTLGA3oq
+uWCEEQejPrgWQyc1tIRt4u+xEIZvHXwFyQRmHAri+b0IZp8hI8ws3XyNBFcc6/P
UZJ42QjYrpePY1LK7yoEGw4yww7Zmij3EeyTtY4dSJqx1jgBTcizLEU1cudLhaAy
55CJKoxE/x5vaeNcvSXVlA896gfVV8Rs8mJrtBBNA4ahdS221Nzl+F0lfVJHw8dm
Il3WpY2gho0rWvNOiQoztkiUa18iFmfm5Syh0zjbAsbF5oQ9f/1oWResrI5thVYQ
Ai5Dzcz8Jv38Se3Lpy1MFhymlxa8exizjk0xm2kR6N+Lu75Re1LRObjqKByYtO17
LAlH+P8ZHjfpuvkxNYOVSVWsGx1/ijW5n1acalOlpPQNTY3TMHQ+Ohv+28FsGUeO
qeC8oVPf0/QjoH/8gDllMz+lncQTX1Exu7wmFzAHD0Q7/VcMOdnxxOLXAYvKgcVc
sd6jMqmdzFIgI0zpQo3kuVlzfIybB4cSgqk7OtQMby1cbv11b0SPeoGeAzQxIXY4
xXXJBxq1yYjeFqXWMA3r1SYXulwxTB/L5m8rWU82mztdf3OI90XCN2Y+b4tiDdmq
XYdAgpYhQYDxXMJhNQLe8psfqzB6Yk/pynZa36/9UHeusPdbEzsvD6LyVsXDwdEB
iBD2Sevb72A1pt2riC32pMz76noYuWrwEduvGQYt3HODKh3o24Uf61snC9AEM5Rz
rzcGcNK3NVPKelFxpz9xzJL3EJyt1uzpFKpgZUlrpkOeli32n7d30fI2aGbIvW7l
iQW4N+NUc5UpcsgwzkE5AIBeMvkk05yvX6N+yFehJKgQlOhtbD3WHEDvHi0VBtEX
NzvL/95UgOPjSYAP73a/IFbtGr23RixUm0mphknPUfNRvWm2D1pksaklJCagIPnN
gV+288eXB+ghWPEu+EZ6RVo8ZG5wcjDRYH7C1Cza3LgNO2q/Iy5VnYkFaelbQdz4
FOavQZuLaAWaBAMfGakq+LVWpKl+K3plEJrb+gLX2iaa/canagWtVcRJVfzB9Gg/
7Tk/Bnin/Q9eHkqL3GRcyyGigjQ5gcNooBCh/mbMLn16Vmhxn6GdGn4Ci3gawNUV
5WVhayX2m30QmSCNjPIDdTG7zufCHp1E/nAaAyG98xeuRhvXu35ufme8dviuR4GS
V7nfPwlS//LV2cl0CAfmz3vcEN8/iisKOzOsKMQ9KhScY/Vt+zKX9xPDj6UwxAbv
vu8p6eS7hH4EHyX/MR2cStxjyzrFho7N4j1J+T9CbJZpV1LyGtMv4MCrG78st8St
ZqkGNyKPJCXMi0804LVMCGIPrk/Cva5/fitjTkwoR3jNnYYbFBOYw2n6DQC8OLGV
yr/MG/MJdgPU9ImRwwZKPbVd15+vjVPGlPFNbSk+zwVZ8/ndtRlf29aDrs2801Jp
VN85hCV66TX/MXDj/kkGtpD41pbZ/cGcJV86AmBnm67bpP67Bo3Dk2en53GmWQpX
CCT4o26nKha4fq39OgVapaKNjW3nJNnvkzxLc/hQURe3meFLi5maAInQlbTOje5z
mDRy8YF40kPdiIXypE5sWwJsxnH/JaMSYgQC+IaWi+estoX0x9heEtrLRa38Rzph
ZiZUZd+rVaiEjwmywVbacUR/LiGWRSENWAQlWeb/ffvUbvHpgLEQkHz+x7qgInqE
LpEyD912hqEVgc0FgvPZ6EuT2P/e81bBWj7XnW+67Ihu05phTNEvFqrYgXg3Q5C1
0GItwK/ko6h1my68ZixcZi2DvuPJAHNvkPiyoDdVS5pdVs3Tztpp6kjWzadhTsbX
3Fro15hLdL35hW6pVYUGnpdkfAuD9eL8mQLYktsVTOubr96+pieSc9ePxcqUyHTC
/BGsrhOSh92bgOeYDKpCyGUedtSedQV2pzWlp84zdw0tY9VmqD/ZUdHA5x8/NrT3
gZiOEtirTLQbUjfEdpLXvNsXHxETpDX2bEBou07XcHLmYtPRHkP3fXMHJD9CrVab
LXE2NsLMQgOqecXlSdqygVU3Qb96zfEsS5EYdhtFwhIAda1ByjkdTfBpT+ACRkbz
dEHG8XXEm/pDAB45wwHiy09rZ6Tcq0kEzNYBLbNshH1TnM1//VrEJfI125BF6+6Z
1/nzXpHLWtFmEBQpCjNU49VMgkV/9gO0hVWi0tFBDbc9qtfd9yeM5fqokc5Mfusj
Z2bFsAvTFeAxgXNz46OGRrAXZT8dD9OKq8Kh9t6975QMDg4UFsQGoB9G8mf95hWG
T7mEMm7EC3p1HDXOzHCjcP0iKni/jMSJfDpG8RpQF7Phx1bshNngfXCqPmASA4Eu
XtJ/gmJSgSbDrPFVEAMWQuQuYZZAHml3g8ED38jdGYk5F201VZ3spV/wOf5BxLIC
6tb4BYM31fdTaSfBPe1nmpyCS9yL4iLPHDqIWhY/IRw0lw2XMhhs5B4UqYYdUCBX
6BHLgUiFaOdOOJkdaEzUpMtqny8jYa1HmMT3k8NDNUNet5sMqZBiCYTU8GjMhOh8
QjJf/0fXqpBy1PHU8cx02XivIjzS12/gkcEhaNR7pVuG147Jot3nzGDzQdKsGdjr
KleQ931ULBex5L4iporQ4VGu/5RIc+p+ofYoY97ny/Ru+QknGM5YdOY9jvMd7EAO
RRKRvvGQqMF4QcI1+WxY9FhWQ9exPEYmITwMP1sR5GMth7HfA8WROOlHtShiMck6
k2imutoBYC1uilbbF0hKyTqkDjwZ5X/X3/sEYuLuLCdAFD3Ot+ZoXPGnh7m6odAM
nl0TbaQN/jT8GaU1wPBXqF4F3HYlyy/AfQBGcqssoOJQVnXs4tBBzWouMGic3zZn
DVN/0FFDNWCkje+whGwjkvVs0jALqXavKiQvG63XiIHMmKQ58otGI0Pc8D23Fqft
UsTarshUhE+sxrZZqKZlOkIaW1/4I0rlfcIy3TyPxVu8IOaKAT0SpauaBMYakk2/
m7u7TUPBo5jZb8/VfIdO2XBxKl+sbfc1yCroHbtsLZlOyY7PGGfXFk1d+PJqj+q+
oDknNqySPJimyl8Gb3+HEyl66XXN6KWUxl3KtumBC5R6vmId3cEAOuvqW8jn5r/h
qmVjI8k5PosWh7d3WZKyW0IuSgJrWB31DznjNv+17GTd0pRJZUukb6zxusUeHrBt
3oFotImiB08h0KxAs+02vze1Z1Hg4ws7NkYMgKoB6UpapPVRbqwpD/WXWVK1TZlg
7e8AMFHrEC6fbrUfQEby8+eU1/4QraGsXOqHpGgsUdq+xVMjSIWgwTvmVgZ/F0Zp
dCoV98TOW6l3BVbeEjWfhUenEBn8tthssOMe3Cs0bwbEw3Aet5/SKCAzHk19FJ6d
3ETRwIafYRvYqBB0Ota3WmXB+iXfRnNKMB25DwG7aDp4uVs4GlSKrmpxtclcRo5o
jYAbfoPMxNbO3QCeEAyaaWACyvVWbO0lKPre4duanYz/5EvB19sTrmvHFzd8n2qB
EqKrMxSwXxx6IiLz2kawxw6MOkglo1HuGJDuB1dgteLVHkQpGqxWyBU6R7Y01LGy
sFyQL+cdKHBzYOA5i670MvSrzyTF3Odb7PbFD6iapE/BtiErtdyc9ot9Vrvz1gvd
crbv3A9ozl5u0bWVsi5gldqES06dv3HG2209NDc4FQA7SQIcbLUif7ouYLwGJjqB
wyqzw1kQG4AWjYQ3vGkVNLP9xSYcuf6MQQcdPCk7EbmM4CF9res9ijkuJ+C7UJQK
oVrTJLM3WvZ2ry+RbE3BjuLkyzjT++62vBNcRAhIQXLPDMdGMurTKPEW3RfpYZTz
ky46+j0LLCyNB5XQN4rDEBLc6pQr3NDodwLhXnDlMFu+/BeATIlkLNWFaRJP8ywU
4D4q4F/YsK4jV7kR6ZSCON3Wo9fOGvoyZv1uZtcexB4LJvLgqR/9QwBz1+5O+MJV
ECo6DraAViwnAqdVCfgOjdpVnTujRjS0Knz4upN39xKiGONJVysYCmMec90J5OL2
yGyFOEFfJ6zNPDKO0NOSMZXLoacHAYnHVTxm9C8T2ysGUnKH+Txuit9duwh5WH7r
SSQ8+5tjV5oWDYOqgQ8hepEScABY06alP5GAhRkmVfOjQQF4IxCml+x3L/isnzOb
pDcsE+CggH7kPIX6eEQirR6s+kELmwILyQZ4dSWuY4EvpjwWVPlMrSSFmJ9yVX4s
xKIgnlDtfS0pj4raw7xByWt8njlDLow1l7Ck2ldMw4erMqJsY5zTWMx3Keo6k5uc
MGxa0hi8GOgddbAhyaSQx6QSEWbmjJcw7dJm0/cHeoNgT26QUOSlM++MHQMmuyUM
Rl5TcnpYOiMLNfau5gM8+X8wd04ivmXk0FYVG/jzQ5LBAwKxwFwDeujTrnMongpt
8NzI/F+n7v0IOFQOqTdRELeL/cLrnn58Z0quUZ5lqZ/VCICulSbtOTjoZ54C0zI7
GzUUU2Vw+r0e4TjhAZT4bKrKKvH+krUnU/7iyHTZ4CRw9/E1jL7y1r1L0R2KY/qO
AmNpXFKO7BiGNlm4OtM6PLymSMU5H/+bVajE84T3LPu2c4Z03/qN6TmClFIBNiI4
86oSc6OpswwijmKjY527VX4sFOY144X6lcJYaW8i1yL74d3APS3ts5f+ZMULxr1D
tFipec84CZTbicnm20pGxLk1imYzygEzWE7tGqt2cGtxUQuAd4ubwXxTUck/G1Jt
BFtNgT4YGUpmtnchxLXs4+ODQsVFSUP6jaCFC9FMK5lxJKV7+fuk7I3uptzXrmHt
R5SjG1+7dvWPcJADhcAajTEDQp1ltdfD79Tifv1zI7Pott9AnZAXIPLuDKc0o5RZ
Gp7iuVSloPWYPnKHm2pedwcAJbRCzGGj8+3DW46QLXHtL8nDldwDrR0zy4jBtske
QVSBgv4l3pOVIolwAWnzzbtZI6Bioqp7d9laf5pXlGStYAzT8ch8/KkPqfyHfMmU
xIs2njJlrwzd/evVD3+UN31eEigyXeVxus91OvUlcsWSWUPX/odciPbV3xdSiQ7T
5QeXAbQdISQDnY0YoUFDMISQTDzsbKEE8lsUawuaLsS7cVxcS9xvSUOT+Ksp/iHp
ZKZ+RXwYpRb1xEcntM8SuZEj4IsIGXwGGc+BkIFCb1ewyQkq35ZhBxaXfsu0Euk2
3D7e7JjJuk8mSK6aAlwlZ/vJBVJ4rj28eN9M5Z8g0s0UezzngVrj4mdQ698FZd0p
W4gg0W8uvYfn4amyaY0qRJUuEXqap7tOnmWPXa24aFPC1DUM0BiCyRqkO3PKXFbc
snRMgCx6OipM8we/x2AV5LW0ON4a26ay1++1V7OwkJRgL7xFuYnqqNGk3apHI9q0
DJof9l/yWmLg4iewmXUp+cbbPjOjO+cMTvE/1c+dYsjU5aia8XwXbg5u463HFicf
2c4mup78ON+aaUcti9tFNZYWZatXKUgC0yZ1laDIHst3AJCSQefuA6PcwWXIBerR
W7QvT7j55rWAmJqLA2AJhzhgP9+dlkwB+CdR9APb5jWs5JCNZWAqzNNNCAqPWVaF
wGrcD5CW8dfUUAaEa0Q3qdrT9dkCJd0aGYUNTLirfzarMrJiOEX3n1wOOrIvPRbt
4/1Y/+TyF+mikL/LNShGPVqxQVbY/DWSwk9IP4u6FsdFwHF2Mz58m9dVMTRVLaS2
TYHGDZx/vUXrMdQTMxU8ZAEn1WCK17oCjQXqrTdNPP6IEnllvpl/cW/ODIHhXsNw
fX+vVwOuqWEdEW6kze1UbFLQ1uTuDD2BXMhO6ILKplWsKJKOzLhXC1aImXibPuQb
8dWFbZGiT1/Tk2UVDYEGp/Up/TaRWVq8c640VA+kC+mCi1MRIWcX/OfPCQkWq3OV
r5UPmxALchhrgGfWpsLm4ncc+AoJan/xXjAZTI2Q6ZIHfIn3Oxg1CwwuMOtHHSgv
S0kUivOoMhViW8jHLlQY2kb7FmjTnLiF1DuaUTAS8P24KOyLARfKh03PkgwqPHz9
MNHJI97lwVCU5zGB2+YQrc630gi8HdiS8p0FKiQtvQqlLxuwQc6J7V5/ZAFHamFw
QLbi/36jETpn/cgq1vvhd90EVozh2jubzumXYQ35T/egNt58MOYOjEFKmNTH1kCU
yYkKpK16ZS7o/27R7UviSeW6Qxp4QHQKNF7QHf/HoaI6M0tYU+/ckpsh1g30zJt5
qMUUKN0o6hT9RcW0MbW7p5CzNcm/maj+B1rfSxzJGtxmEcbbq2mnukYm8yVxBBHS
hrQk017/muXpf/IAWDDOJUWu6Fx8nVGH3hDyNUrEk4WCzgYIX4Je1a3I6W3I+J1q
wghqI7YyIuW0RVgEmln1943DhPWCiA17aM70UPs0NjXQALNxQq/Whee/sBrRnfjO
Ae/0Ps5iEb3UWb8XU0KyHijoawHpS6XeiikeETe6wUZwU10Q/XeOkhNKVFiicBrs
YNrVbRXhUBn7uis+B5i9XP9AYOLdPlEcHkxom68ZdRV6K3QtgZuw95raGlWpFioS
JdIIgp9ffzoqgL2hRMPXx3H5krwEK6fHDB2St1M/+3T8cF2ahl87tppLStG9Nf25
QG+7GA+S22SEdsdjKvi3ggQ/vp9Y08lFMidcXMFo055ct3+rZASnSjkS9ipbkPwS
tWvgyretGmi7uFOmFSenORzHt9PzqT8cxa9iTFo1I9XqO1Ec/pekjGI8mqHgUK07
QDnE3NHzhtZcLNNOEAS3gnmZzVvmpKlpw/k7r3fyw2q3/T6xvbLDTGb5V5OOsOs2
x+y2035Tp2JirYw4TYEeONsar5zljwHzHcy1pnAzG4njNbiC7MYACG2zCbEGtcTG
edntACC4dIRMQCcLyhLHklqZDzvwJH5IkS+owFGI8BRRU0brknWXfMgQlQrTSC0V
9pYCItvzlNvohguWucJ4iKTQpQwxZ4zN15I2QjuIU+ERKaL29SxZj1BP+LVFrdSp
wA1VFSaekWjb9cu6+cpsW5bXB5E1qZ9aC7PUrJyyZV2cJQzsMmyGHhyNasVrHGG6
slI9NZuXL+//HltHu8P4pKdMpIZab92x42KINrnufbwDBZy3GfNWno9JZM3xBqef
uytOdmpVRRMPByDC+DC5wWFTo9CiqSxzHvAqdzllW0HdbFBVTC6n2/EYZzq0Stt6
C9pWo3qh7wAe+AmyfIsIETdMrEvqUswek4Nbxv1W0lU0X2GKL0e9GUo0FvvD8PvP
NJ3a9e+z4ODst5PvlAP2nXqMPEsnug54g4+AnOrQN3T1T1p7BEAplJDpPOUzLciM
MF1jmM5eE3XUOPJJHwgE/aX1D1P3lkNFyeKWkBnRTRI6MEl9fgVZF2806lYpNe5Z
Y8H66kjy8oFBUNiRjuB4eeW8gVqDkpB5cRH5pnxGSGURBRNcWmVBPnj5Lvfh0e0u
RIdRlx2DMai3wwPl0DVSDQNqbaPGN3Tx0u6RWeF1OfdZCJo1GsKqXQH9X9Mm/o0P
dhwmYhgh2jYL1IC4pGHqQw5dcIXMsI6EHkFGh3exJ5X7zvOHC+qKkEQhUOXypOYX
Kg+YxpZ6d9OTcjHGywBuKThjUHgw6+GSmcjRi+Sphb2xaVoXhQ+NZeom/lslOIPB
9f/Af6uMgxCfKmiyUm3GsPT957YUujYz+eVW6aHrFQgLWHGnT3674qeoL9VM/VrP
cHG5m7OiMYrnVSASuBSBw7GxYVtcxejO316/05UvfOqe7KvgRKdyxDgmUUFj+NqJ
sIosUp/3S1saQnSSJwq99/K3Tpk2TmmuDdmIzjxAynMXT2wpeh0qPf3JgKzDZ6id
K8JcgMSV4NejkPNfmrvklwdMNa/5OcGCAPzp661vgn7UniKR2WdqMy4kC84rkWKv
097qFiFT63HmmxN1OsNdyISRn8oQwhlH5eWjtyjPy2rM6vvfj3SuRgLhL07cE70v
ydspJnG8IhXJ2w779P6zlvqFqkcmNxvfqtwEh83on311wD3D+Z9z9FiHbw3aanHV
+Nzk/RvlPZ2s0q7lo7rs8uo1jribDjDK9WtPQ16zxAT4F/Ep9Z27TexkNIBUSQ8h
R1qGIlaExR86ndr76c5LFTRXMlfGl5ICMi9NUcDRBrHFsecw3Rqujjc1EwVLVk0X
lVY7heI8s8rk5ompswdIGrX64Ms2W2KV81XEhmyT1HyFh/MVxdss9t7IODN8H2Kr
Lnr5JWqd9xZbTuMcxvxjbhmzFUtTHnGe/+fkV5L3TfGE70NTckEn/lj72gifbP4e
ZbilzPIRiroYWuJBdhmJ28vBwMmpqZMLtKZg2qS96nbfKSvqbbW2xQ+JyK8+Z4/0
yf/J/0XP7P4V9OCUkYQ/qFyd2QpUylb0kL5GWsDrSoFwyYjO3oeW0r41DPEt6WRv
VZmjETfS7toftG0KSCeFJorSGBd9GWkEux4GT4BR3XjE6V+C6bwXiwmWFc9I9Fkd
hddUIerNeNMi4g0h32lfw70zEAxKHSeMSVZKk99HDw9E9+GPqsJgilLYzS4WKQAs
CIFlPMIMw3z016xjck14pIJ4n80WVLbeSG56+/IVFZ5PIvlBZPo/mX0eYvj7Wo+t
Tmrewe3UPIUNIojn3u+ILL3xRSz+1Seli/I9S6dJh704r7u4Q0HEHNmEo7GFIDW3
38zLfNKG0XTIJI1QdPwsZGCTlA1iB7Tgx3rvsKcrJyiAXw+irDQ4wxGz9Zmd6wJV
YH2CESWZ5Yz4Z/0OY5DznrpbkNQEPh8qAx9ptSjrsv0OuLrG1bWNzzvE7OLnDkUH
IHi7Jz14Fhui36RBNypTvyqk4Fb4r1GAvbdHEsabdUNS7LmntrRLpcZs2a8d272m
KurT5ArBKu8N57Y0/Tu5c6thcpzGFGaEzITdnfftYzyGxsyoAfnMf445szm87hMT
DUwVYiXhYBjBZiKWMa/dzgpHb65JkITGIFHpXDCaP5DTiTpImwKMFWRPVY61J6mM
2cANFSKTkGWF8FHF8htn6T5JZZsquxXmU2ssOg+2pnqVy4FfvpMvB1bbeDf7Q0sg
BHV0GvN/cOx5kJvGkG/mTlvq2hu6jP9aYlKYbE0mHYOayCCFnSY/f91ND389Djau
LnIvPfmiVSI4OtHrRhEuvLo2xWcxTDISsEoe0c8AIKSRFn1uM7cXx8zt803RPDHx
ZBPMhvjOgzBjSCic5LcqQN40vLdxjbdwD0L6k4TfJT/jkvtAQCzRfRy4KY523eA6
U277TmuDq3G6BISRlZGj04HCtrmq0zHPSWnHwGN9NHp/vqAo31e48irSA1xcL3gD
fdSLhHOoR7/gR79cWWWD7z6a1WeTWliGPaCELhhb+XgmPKOHjRSEajS/SszviQGl
7xWxbciyjpTEIWKBaTXWRpyYVFldG3muKKMkMjDh10md7ODagqWHETuAg4UWWo/t
7a1lpZ8mCjdmYIpK0d96wLJMwSefKxtFut1JKQh/gi1LzwpVqStcLizAOgB8VHup
YcqjqQ9Geh0lxHYceLIEgOADENK7ACmz3TZ2nQa0hNqi0Vb3/kwl7da2SNj+XD+v
IAmknr2fdOhXr1vHbqEbnV8d8nhokwoyTB/gjlThA+8DSsgXZusINIRRw/tA+xg1
mm+1gGTEyKTujFVaC7oMCoB18FFS45Xzyw6YSkFsynKLhfoK/+Y0uQCXWnxqYQUp
i+giuNSrucduX4r5dYNwz8Cf5SYlsNYEWoDQNFm8npFl/l5YjmSudDGYFvCvBCWA
DAC7M2/oo0/uA1jLR32ZKPpGktVy4dWT2N47rY5FqzfN04N3O7AbZMMTIxjI6tR8
7gRWqiVUIImr41f9jEqi6wDlVOkJMiklCvjXEzOebf5uQBZqhWaDWZAVvCdhtMk+
em94+whEF/IDo2hBB1AO7RMKUp6DDsMSLE/koA+dk8+Vm+LSuifzzox8C+vAf+l9
lZdzVw036jIC8y5y6AX6XJKH2n2h0rWcu1QU0UA5QTcyPCod58OGJUIxcT4jCOZZ
Fchti17/RiiC6xPu31eWUyyBKO/tjHAekwoLvKKKAjDzzsridg8KJgq+THX7y0Bd
lLUtX9p1AW0R6/USsc0bbObtzIlPmOBDYS2wWkece/3uN5biEU/9APpgTUEbsqk+
F++qsqztuw/XkRpn7avg6SiE2CB2I6vEvA7C/NAgdNFIGk0mchyXaNZnTG6Lb+I4
ydY0Y+qOYZjU19skyq8qQ+l6bL2wIOyMlDeZX5hIEfLvXyZNBYjiZMhaWYutccc4
v8FlDKuOZju4bmQ02+aLAmSRbNSwKhXxQu4AP6tXenZaHntYLDOty+TxqgiL0fJg
ivodg7iA2bZH/RUe7c7OZ++DL9OauSlkjhnkKfcj+vWIFmvE8H6sl5xJ8gjZoS8K
nEVq4APspjcXmSu0JaqAMyivKG/cMkgSa9zM4U7Nms5GkKOajw8iA1I6Elri7uYX
oBkBBJ+BhK1wvoC+L6UKSGSCuuLB1zZM/SeXlNRNwRKViuC7Zh6Rl0/1ejpJ7jdr
T/eEbXkz1yae2IKRFiHO6xQxPvRiMzv+U7r0+0+JHHUbtNDFPYYMHeTNyCLbhDXC
Kug+pTjj8An1JuUCuL3CzqQXsvfD3wVLteFJn3NYq39XtFRLjzBT+mXYsxQv0hnr
5Yu2py0zQ4Bh2NoLidT8VQTA3I6A+4Q/gtIdDa/omb1xyi00pAzt0kOemWRxs1o0
y27oGetSX1UTYnXp2832JBV4xq3zQEBLqbRIeY5mtzt1VcjXKJkBZU5oaDhqHe6W
gUXvB35JggEXOxpc9sOlpser9KrUY7MTV+mpkK1/9lPfda2tcbiDjBxWnoZK3VKa
SQJpzYy1WpdilhLqe1aOwgNBv7So9G1ThuPLFv5OFRwulxEoCz/Yw7lbPZH0jKO+
oFYFrsIyM2gvR63vZH+sDy5mgHriXDxjQVtCz0+PPxEWfdFmKTjCFP6lRVxPjWKo
3Xf6XNfqWuLUdy6N7AHTnzjkW1unkcUXkES47f/Rf1w+0xyzdwb2IELlKuCtZj6g
8aa84tQNyNQYgjZlygpSv/4BLK1Z1vMOB6eNW3LKkYyRa5XXk2wtOSOTnxurELS7
fXir4iGHheIDj/WpRXSrHba/mr91n3S25dDhFUcildRCwTSztHtZry2J9880m/5i
cgH7kUhNW2/jfkT1ZA+ePXRQMXa/+DCwAJNY3Suy4J80mp2hQ+5MrRHiWHKiwZNO
1YG36TxukXFtsVsCvlJ9tWE2DxXjr8Qbgnk2nYR/0lCHFpW7yX6dKq2Vv7KSTlK7
k3P4AXU/2Q8qztqptZbME0dWwHJ5ldB7T2WvMEUpIzs93HhbgDNwOpfPFhpvC09S
vO8hot1UKC2ZmHJsl6s4kTFFa9z5YfJoK15bHjys5piZ5r5h83yYADwvOGD0BXEa
YAvOTHShkz1uGAqnBzJxKoqSPZY3a5GrsDsdD4JF0gK41g/za8kfF1/iyrZCQ9I8
WAbgMA7/hPCN+sQp+MOPxh8XwYEvOQtabO3z6BG1+jDHGdcaAtIr9sq1Ccul/+zb
nPjB0xYt6uu+tFOlHtvxKmXEcNPOUifaMX7rZPBUwAHemgdAW8dRMTxVnV1zwNVw
C2sSY5VAoDaESkDJgQD0iQQoqPeol1+U8hYtJoQ/1vS/IlztlsRmqmMbuT5BGeQt
P3uxbeYro6jgEAkaurH/IuoKANVDUBXvq2srpcM/TDD0VksedIzN3AgPSw++oaO5
MQ2R1++8QkoU4mBmjsVTgDyM/ifDDQjRWp0W4nl1GeyL6Rr4y4akQB9SNeHdRMvq
czZXdX6Jv324oFXMQOzXQBsWCW1ro36Aw6S5WIx+xkg1sEqZlgFE4or8CAFX8v54
mD8LHC1I057/OjyjPGr3b2I6hBYUUbrx1mqcrH9UEP46HPlZEew0R1InPsW7Ewns
41pIgNzXy5/zoUIM/yLj76uPKmI0Ea4hOMu4IY9RShFoMgQsvEGQlwrqv+lYerBo
21uPBqt4p1JAK7xPlw+aaS9NAU2lCTNfsSVT2yVIdnHce1Ih9Pj9QvVH0EkVjMSP
jSoiQh9KhWMe/CdbFQPP0/euSxERujBzwy//2lM5hWxov1rnBG3+479wj8rBf95a
k/86AQHBQRwEONMVAFDv7dAPSzjfRIpqpM1RnOzQBz1U9H1n/qZpuasYHAUvs7WG
mMqc9RzHCOrLEu8O6fhbuUVTfH+9bKWpb9oieW62rEmOvObEDuVNxTfg0JQoGpXw
f0Lhb2/II6pC+r0fz8sBMmN2c0aL3+hSRQMH57Akw2W980K+0krIzGFBQ+X87KIR
0yTHCT9qn3iH2jtzRtVh+Ynq7YwfEr78OVFx87hDOErIkOZdDFfT6MTbZQAMp1LV
bp9kYpRA+QInoGqoockVFELcDgbn7htFI3Yr9Fhhg3+StdDD1Bd/4BwoO3mI9Ogp
j6I1Ltt2E88nCM/7zuNxyn2RnKBryoVAdfwHbfih/9nZgO0upSml/PC8NTQrMXJK
ju09Zc9sgX2PIHtyVAniMlxZqyIGiRK2zo5ljWVzdeRNWgpOEtIbckEsPf3GSjTL
7ULMDvIk+TV0KttGQjFguYo2Gn5CgnC2o4XvVpty1p+asExzjVGIAa9ia/Sermup
+c4TnYuMRdzDEk+XmTJchThWwx3+uaTeQ+oCebReqUVHSuqvFsAjpZi7VNz4OvQV
MkbYn33fvuAndkHbjiUcnhJOPhS/RxuTJtmMu7EoBnXHm+Jouu7VGzdhgPzQXGy2
UBNJJeqokGDWcn6jTYnBK1YCgZGYOBBF37HLwaSpYqknJhK/cYKx9CxIYJQVmmyo
Ed1nYACkUpiObRa5S4wzpcUk4jwbjdIVAZodmUfrZ0RnABZP4GsYGGaG1SUmHYQz
t8iTIatZWQHNkTF+JgTdYXb3zzK4DMKL4ocURNzSCUOJB+h2iIi+AYoGpJZWa6FT
O+pQJAHOJcpkz+Cf/PXOxUANAT4p8j4C7JD4s5uvbDYAyWBC7vQsKjpwJAycBo7H
lb0WMHdcKfUv86R6N05N5JkaIdzbZ0ejfBIRUQKUN4tnrvhL+qldQelVnUKhTiyL
Z1FUEZrKTaGy42XF54ldloOoRDe/Lp07imiXPZWjgjbkvC45YzC48qIyKDE6Z50C
pysta9tNaA7SAj5qMOQtc87vtghjdKqU3v2xwRywn7HZr+IZFrTDZz3HzLGc4tzU
1dQ5Mq12F/YgwQaqKXCLYIdOZIOovz4LPCw0BZ7ohlGqQQMg98c2g8OmZfp1G6sQ
2+HUDcHJpSXDQ1o+phhNvDU8fIiS2OsxqiyQmmoLgUtubJqbXzzy264pm7kvAJG9
oWxOfbp7XSxLFo7R779o8l6XLuoYsP2uud1GjG6E49VEIys8QVt18tUFfwq0n43t
kRuIqh+14NkQD+3oj23DPlrkF94aWgQp8RUDyAQhdaG3Pv0meFT2NrTdssU1Kd5n
tOYd0ybag5J7v1K2sVLLBdHezk4PRpuiwzBZsWPltG+FpaFyGLtOg1wrQtMC93Ak
6dvRwVKWLMmA6KCTgqcLSZMhctZyfDGGDwaVBT3KB9GybGQUF+yc0+yjlPZzLFqK
PTf34RxgDRKG1vf5HihxShxYCQ88/MDEDv1tRmy0Bq0uZ/+WPZzC7OcotdenkDxF
fvjDz8l6/F8PutyL3Zs0lzTvzac5vGNAq36i1YWiGNeQ+QZGxQRCspZ1D8BITuXb
BJqAmFIBPlMwoPTj2mrok0v3iLjB5iKr7bHA8XByTu862rs2MTQMm9D7lFDALne7
OjL2JIWq9kKYMRq9UjGwZNV3s8PrMWDrIhNqVmAm7B4l2yEJp306Gc2KOnOBUfrl
egEDsX0jENTGuhVz3iVegEI8h7g/HGtueln2NwC8Zcms3eiXHi9baDpv8hrhREvW
bUkcGbmf1LOSFkC+Xqi2lmD9c2sJFR8BPNtxX9YGS/oK7OlC6uK7Ad2V6KKJnEHX
6XPQDhI/jP0oZbBDKm2+dlivihKJMy6BNtvzod26x9Xji+15AotjqON8hT4AgoG/
uqpRWBnlKBdOnTx36VaEde265PpAsa80A+5wlwC9ErKb4cHl406bOVdRtMfDO2xo
HCErvaBgWmuaxk+F7E5xkL9CzVnCnQv+k1XeRwDTa+qkIwD5LQ4b8gLPlwZbBysw
s7vzrMb+NouPDbhMP1/QiGHXTb8ie0Ql2JGZo8dgxj7sbu4jZ85ntFj0DxaFPTEi
GNrKJ+ac5Nc9vbLSi0h3PyXkdtCYUlSE5Ix6shdrWtDy7nR36WlRDHziZ/XeSjW4
0qOJipeKwRc5FX/t0dLh7uPJyl/93YY8nAYlHmi5JE0FYUetZtFnu8FzvLnIVIYy
BPU/TYoBLhwlfX/UC0Qg2YvO+dqdTaOKconEremgn+HlOZqCDqLnsXhKSaEFqVQX
5kZFrDLmMKUsfbLVy3NbO30Ny3DFjkoYB1wgSzU7Yr+o7IcZzzdrFrtmPkhwE+P/
SiXXmicgRrbkoXhmqQnIBlcua3QL902chK5IRvW0DM90KW6V96mI+t4Rlyk5CVKS
ZySoi9WUMQSko3N6PM3oQ2dLWA1btz8r0GNS32kcPFhRE2duEpA2Sa0bR3jIDep3
fpkd1AJyaXluh4UoURCtbqxRHIsSs0x/0xLqJM3M3JaFG338SnAOwDaAlCZlcH2e
Nkkjg7bHab+zOtqgbMSwngERtA9M/MMK7KjzlBMLf5Rbb8IfkfuyGNnCX1ifEaTt
psRJ6yj3N7nLzsKNMXxR362TaY4cx0umIK8eOmLslyRBgY54Oi3inhAsaq45Z/Od
VhlcvPqjGfhz+JGWYMMUlwzGf+XwS6zEr0g1uLr5gx/y74gVfxxOkB4YbdTjGWrd
qT3sRv3lR83mw6dHIBGHgRxvE95mf0f4GubMYS5yI+E63Vhabpvmwvws7WgjibVY
g8R8hGLh22J+g4e8j06pTGMVTWe6SLH4YbrBbaw22CG7ovcsutYnlq+y76XLcFAE
63QTFgxIupz/iZd5phqrdTUkX+/ZGx59dsJ6dAoadZrJRktwJn/X2VgxhdgLHi9z
TCAAGtvGptM5qQkHJQlEaYhFqBo4R4GVHyBZa1c1dA0klC3xZDpcZA3yF+Ii+uEv
pPKcckkVOZbA074TpLllj5sdxXkxMZA806rrRPZWeM2x3o9glUK/IwD3tJ11OD9S
rCJF0N9CU9p4G/+gJ93lyV1vRo5SLG8JynQjK1V3d166ozz5Dozu8n3S4vSt8U8U
yMfaUmEs8HgdaX5z5wgfjVPESwN3oFWycuTrR6JDbCQB4mULFfDTyvymC1FY6kXV
VxWQGhLrVqgga+4/bcsHfCOc7pH8hV7sdh861kT/YDNLzyQIzjZ3AQryLjq9yD6w
mwz0YQE8XRqiYEoh4ZkReTpDG3K1GuLW6Mm7ZEDiGLArmebayxQjO4ED6oUV4SyN
4KbvBksnb2aOvKrwi8UJJThrHsCoklM0lz6flxWEbVfuLsQcFmrFP7mOJxHWRESc
8ZfiJsTZ9LleZaf6nFO0eg==
`pragma protect end_protected
