-- TEDv3_architecture.vhd

-- Generated using ACDS version 14.1 190 at 2015.03.30.18:27:41

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TEDv3_architecture is
	port (
		black_interface_mac_mdio_connection_mdc           : out   std_logic;                                        --         black_interface_mac_mdio_connection.mdc
		black_interface_mac_mdio_connection_mdio_in       : in    std_logic                     := '0';             --                                            .mdio_in
		black_interface_mac_mdio_connection_mdio_out      : out   std_logic;                                        --                                            .mdio_out
		black_interface_mac_mdio_connection_mdio_oen      : out   std_logic;                                        --                                            .mdio_oen
		black_interface_mac_misc_connection_xon_gen       : in    std_logic                     := '0';             --         black_interface_mac_misc_connection.xon_gen
		black_interface_mac_misc_connection_xoff_gen      : in    std_logic                     := '0';             --                                            .xoff_gen
		black_interface_mac_misc_connection_ff_tx_crc_fwd : in    std_logic                     := '0';             --                                            .ff_tx_crc_fwd
		black_interface_mac_misc_connection_ff_tx_septy   : out   std_logic;                                        --                                            .ff_tx_septy
		black_interface_mac_misc_connection_tx_ff_uflow   : out   std_logic;                                        --                                            .tx_ff_uflow
		black_interface_mac_misc_connection_ff_tx_a_full  : out   std_logic;                                        --                                            .ff_tx_a_full
		black_interface_mac_misc_connection_ff_tx_a_empty : out   std_logic;                                        --                                            .ff_tx_a_empty
		black_interface_mac_misc_connection_rx_err_stat   : out   std_logic_vector(17 downto 0);                    --                                            .rx_err_stat
		black_interface_mac_misc_connection_rx_frm_type   : out   std_logic_vector(3 downto 0);                     --                                            .rx_frm_type
		black_interface_mac_misc_connection_ff_rx_dsav    : out   std_logic;                                        --                                            .ff_rx_dsav
		black_interface_mac_misc_connection_ff_rx_a_full  : out   std_logic;                                        --                                            .ff_rx_a_full
		black_interface_mac_misc_connection_ff_rx_a_empty : out   std_logic;                                        --                                            .ff_rx_a_empty
		black_interface_mac_rgmii_connection_rgmii_in     : in    std_logic_vector(3 downto 0)  := (others => '0'); --        black_interface_mac_rgmii_connection.rgmii_in
		black_interface_mac_rgmii_connection_rgmii_out    : out   std_logic_vector(3 downto 0);                     --                                            .rgmii_out
		black_interface_mac_rgmii_connection_rx_control   : in    std_logic                     := '0';             --                                            .rx_control
		black_interface_mac_rgmii_connection_tx_control   : out   std_logic;                                        --                                            .tx_control
		black_interface_mac_status_connection_set_10      : in    std_logic                     := '0';             --       black_interface_mac_status_connection.set_10
		black_interface_mac_status_connection_set_1000    : in    std_logic                     := '0';             --                                            .set_1000
		black_interface_mac_status_connection_eth_mode    : out   std_logic;                                        --                                            .eth_mode
		black_interface_mac_status_connection_ena_10      : out   std_logic;                                        --                                            .ena_10
		black_interface_pcs_mac_rx_clock_connection_clk   : in    std_logic                     := '0';             -- black_interface_pcs_mac_rx_clock_connection.clk
		black_interface_pcs_mac_tx_clock_connection_clk   : in    std_logic                     := '0';             -- black_interface_pcs_mac_tx_clock_connection.clk
		clk_clk                                           : in    std_logic                     := '0';             --                                         clk.clk
		hex_conduit_hex_conduit                           : out   std_logic_vector(31 downto 0);                    --                                 hex_conduit.hex_conduit
		input_port_external_connection_export             : in    std_logic_vector(31 downto 0) := (others => '0'); --              input_port_external_connection.export
		lcd_clk_areset_conduit_export                     : in    std_logic                     := '0';             --                      lcd_clk_areset_conduit.export
		lcd_clk_locked_conduit_export                     : out   std_logic;                                        --                      lcd_clk_locked_conduit.export
		lcd_clk_phasedone_conduit_export                  : out   std_logic;                                        --                   lcd_clk_phasedone_conduit.export
		lcd_external_interface_DATA                       : inout std_logic_vector(7 downto 0)  := (others => '0'); --                      lcd_external_interface.DATA
		lcd_external_interface_ON                         : out   std_logic;                                        --                                            .ON
		lcd_external_interface_BLON                       : out   std_logic;                                        --                                            .BLON
		lcd_external_interface_EN                         : out   std_logic;                                        --                                            .EN
		lcd_external_interface_RS                         : out   std_logic;                                        --                                            .RS
		lcd_external_interface_RW                         : out   std_logic;                                        --                                            .RW
		output_port_external_connection_export            : out   std_logic_vector(31 downto 0);                    --             output_port_external_connection.export
		red_interface_mac_mdio_connection_mdc             : out   std_logic;                                        --           red_interface_mac_mdio_connection.mdc
		red_interface_mac_mdio_connection_mdio_in         : in    std_logic                     := '0';             --                                            .mdio_in
		red_interface_mac_mdio_connection_mdio_out        : out   std_logic;                                        --                                            .mdio_out
		red_interface_mac_mdio_connection_mdio_oen        : out   std_logic;                                        --                                            .mdio_oen
		red_interface_mac_misc_connection_xon_gen         : in    std_logic                     := '0';             --           red_interface_mac_misc_connection.xon_gen
		red_interface_mac_misc_connection_xoff_gen        : in    std_logic                     := '0';             --                                            .xoff_gen
		red_interface_mac_misc_connection_ff_tx_crc_fwd   : in    std_logic                     := '0';             --                                            .ff_tx_crc_fwd
		red_interface_mac_misc_connection_ff_tx_septy     : out   std_logic;                                        --                                            .ff_tx_septy
		red_interface_mac_misc_connection_tx_ff_uflow     : out   std_logic;                                        --                                            .tx_ff_uflow
		red_interface_mac_misc_connection_ff_tx_a_full    : out   std_logic;                                        --                                            .ff_tx_a_full
		red_interface_mac_misc_connection_ff_tx_a_empty   : out   std_logic;                                        --                                            .ff_tx_a_empty
		red_interface_mac_misc_connection_rx_err_stat     : out   std_logic_vector(17 downto 0);                    --                                            .rx_err_stat
		red_interface_mac_misc_connection_rx_frm_type     : out   std_logic_vector(3 downto 0);                     --                                            .rx_frm_type
		red_interface_mac_misc_connection_ff_rx_dsav      : out   std_logic;                                        --                                            .ff_rx_dsav
		red_interface_mac_misc_connection_ff_rx_a_full    : out   std_logic;                                        --                                            .ff_rx_a_full
		red_interface_mac_misc_connection_ff_rx_a_empty   : out   std_logic;                                        --                                            .ff_rx_a_empty
		red_interface_mac_rgmii_connection_rgmii_in       : in    std_logic_vector(3 downto 0)  := (others => '0'); --          red_interface_mac_rgmii_connection.rgmii_in
		red_interface_mac_rgmii_connection_rgmii_out      : out   std_logic_vector(3 downto 0);                     --                                            .rgmii_out
		red_interface_mac_rgmii_connection_rx_control     : in    std_logic                     := '0';             --                                            .rx_control
		red_interface_mac_rgmii_connection_tx_control     : out   std_logic;                                        --                                            .tx_control
		red_interface_mac_status_connection_set_10        : in    std_logic                     := '0';             --         red_interface_mac_status_connection.set_10
		red_interface_mac_status_connection_set_1000      : in    std_logic                     := '0';             --                                            .set_1000
		red_interface_mac_status_connection_eth_mode      : out   std_logic;                                        --                                            .eth_mode
		red_interface_mac_status_connection_ena_10        : out   std_logic;                                        --                                            .ena_10
		red_interface_pcs_mac_rx_clock_connection_clk     : in    std_logic                     := '0';             --   red_interface_pcs_mac_rx_clock_connection.clk
		red_interface_pcs_mac_tx_clock_connection_clk     : in    std_logic                     := '0';             --   red_interface_pcs_mac_tx_clock_connection.clk
		reset_reset_n                                     : in    std_logic                     := '0'              --                                       reset.reset_n
	);
end entity TEDv3_architecture;

architecture rtl of TEDv3_architecture is
	component TEDv3_architecture_black_interface is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			xon_gen       : in  std_logic                     := 'X';             -- xon_gen
			xoff_gen      : in  std_logic                     := 'X';             -- xoff_gen
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component TEDv3_architecture_black_interface;

	component TEDv3_architecture_black_rx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			in_startofpacket              : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket                : in  std_logic                     := 'X';             -- endofpacket
			in_data                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid                      : in  std_logic                     := 'X';             -- valid
			in_ready                      : out std_logic;                                        -- ready
			in_empty                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component TEDv3_architecture_black_rx;

	component TEDv3_architecture_black_to_red_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component TEDv3_architecture_black_to_red_memory;

	component TEDv3_architecture_black_tx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(31 downto 0);                    -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic;                                        -- startofpacket
			out_empty                     : out std_logic_vector(1 downto 0)                      -- empty
		);
	end component TEDv3_architecture_black_tx;

	component TEDv3_architecture_descriptor_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component TEDv3_architecture_descriptor_mem;

	component TEDv3_architecture_heap_stack is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component TEDv3_architecture_heap_stack;

	component reg32_avalon_interface is
		port (
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			chipselect : in  std_logic                     := 'X';             -- chipselect
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			clock      : in  std_logic                     := 'X';             -- clk
			resetn     : in  std_logic                     := 'X';             -- reset_n
			Q_export   : out std_logic_vector(31 downto 0)                     -- hex_conduit
		);
	end component reg32_avalon_interface;

	component TEDv3_architecture_input_port is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component TEDv3_architecture_input_port;

	component TEDv3_architecture_instruction_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component TEDv3_architecture_instruction_memory;

	component TEDv3_architecture_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component TEDv3_architecture_jtag_uart;

	component TEDv3_architecture_lcd is
		port (
			clk         : in    std_logic                    := 'X';             -- clk
			reset       : in    std_logic                    := 'X';             -- reset
			address     : in    std_logic                    := 'X';             -- address
			chipselect  : in    std_logic                    := 'X';             -- chipselect
			read        : in    std_logic                    := 'X';             -- read
			write       : in    std_logic                    := 'X';             -- write
			writedata   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(7 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                       -- waitrequest
			LCD_DATA    : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_ON      : out   std_logic;                                       -- export
			LCD_BLON    : out   std_logic;                                       -- export
			LCD_EN      : out   std_logic;                                       -- export
			LCD_RS      : out   std_logic;                                       -- export
			LCD_RW      : out   std_logic                                        -- export
		);
	end component TEDv3_architecture_lcd;

	component TEDv3_architecture_lcd_clk is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component TEDv3_architecture_lcd_clk;

	component TEDv3_architecture_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(20 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component TEDv3_architecture_nios2_qsys_0;

	component TEDv3_architecture_output_port is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component TEDv3_architecture_output_port;

	component TEDv3_architecture_red_to_black_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component TEDv3_architecture_red_to_black_memory;

	component TEDv3_architecture_system_id is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component TEDv3_architecture_system_id;

	component TEDv3_architecture_system_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component TEDv3_architecture_system_timer;

	component ted_crypto is
		port (
			csi_clock_clk                : in  std_logic                     := 'X';             -- clk
			csi_clock_reset              : in  std_logic                     := 'X';             -- reset
			avm_read_master_read         : out std_logic;                                        -- read
			avm_read_master_address      : out std_logic_vector(31 downto 0);                    -- address
			avm_read_master_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_read_master_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			avm_write_master_write       : out std_logic;                                        -- write
			avm_write_master_address     : out std_logic_vector(31 downto 0);                    -- address
			avm_write_master_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			avm_write_master_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			avs_csr_address              : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avs_csr_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			avs_csr_write                : in  std_logic                     := 'X';             -- write
			avs_csr_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component ted_crypto;

	component TEDv3_architecture_mm_interconnect_0 is
		port (
			lcd_clk_c0_clk                                   : in  std_logic                     := 'X';             -- clk
			sys_clk_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			lcd_reset_reset_bridge_in_reset_reset            : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			black_rx_descriptor_read_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			black_rx_descriptor_read_waitrequest             : out std_logic;                                        -- waitrequest
			black_rx_descriptor_read_read                    : in  std_logic                     := 'X';             -- read
			black_rx_descriptor_read_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			black_rx_descriptor_read_readdatavalid           : out std_logic;                                        -- readdatavalid
			black_rx_descriptor_write_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			black_rx_descriptor_write_waitrequest            : out std_logic;                                        -- waitrequest
			black_rx_descriptor_write_write                  : in  std_logic                     := 'X';             -- write
			black_rx_descriptor_write_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			black_rx_m_write_address                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			black_rx_m_write_waitrequest                     : out std_logic;                                        -- waitrequest
			black_rx_m_write_byteenable                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			black_rx_m_write_write                           : in  std_logic                     := 'X';             -- write
			black_rx_m_write_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			black_tx_descriptor_read_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			black_tx_descriptor_read_waitrequest             : out std_logic;                                        -- waitrequest
			black_tx_descriptor_read_read                    : in  std_logic                     := 'X';             -- read
			black_tx_descriptor_read_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			black_tx_descriptor_read_readdatavalid           : out std_logic;                                        -- readdatavalid
			black_tx_descriptor_write_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			black_tx_descriptor_write_waitrequest            : out std_logic;                                        -- waitrequest
			black_tx_descriptor_write_write                  : in  std_logic                     := 'X';             -- write
			black_tx_descriptor_write_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			black_tx_m_read_address                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			black_tx_m_read_waitrequest                      : out std_logic;                                        -- waitrequest
			black_tx_m_read_read                             : in  std_logic                     := 'X';             -- read
			black_tx_m_read_readdata                         : out std_logic_vector(31 downto 0);                    -- readdata
			black_tx_m_read_readdatavalid                    : out std_logic;                                        -- readdatavalid
			nios2_qsys_0_data_master_address                 : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_qsys_0_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_0_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_qsys_0_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_0_instruction_master_address          : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_qsys_0_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			red_rx_descriptor_read_address                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			red_rx_descriptor_read_waitrequest               : out std_logic;                                        -- waitrequest
			red_rx_descriptor_read_read                      : in  std_logic                     := 'X';             -- read
			red_rx_descriptor_read_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			red_rx_descriptor_read_readdatavalid             : out std_logic;                                        -- readdatavalid
			red_rx_descriptor_write_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			red_rx_descriptor_write_waitrequest              : out std_logic;                                        -- waitrequest
			red_rx_descriptor_write_write                    : in  std_logic                     := 'X';             -- write
			red_rx_descriptor_write_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			red_rx_m_write_address                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			red_rx_m_write_waitrequest                       : out std_logic;                                        -- waitrequest
			red_rx_m_write_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			red_rx_m_write_write                             : in  std_logic                     := 'X';             -- write
			red_rx_m_write_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			red_tx_descriptor_read_address                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			red_tx_descriptor_read_waitrequest               : out std_logic;                                        -- waitrequest
			red_tx_descriptor_read_read                      : in  std_logic                     := 'X';             -- read
			red_tx_descriptor_read_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			red_tx_descriptor_read_readdatavalid             : out std_logic;                                        -- readdatavalid
			red_tx_descriptor_write_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			red_tx_descriptor_write_waitrequest              : out std_logic;                                        -- waitrequest
			red_tx_descriptor_write_write                    : in  std_logic                     := 'X';             -- write
			red_tx_descriptor_write_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			red_tx_m_read_address                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			red_tx_m_read_waitrequest                        : out std_logic;                                        -- waitrequest
			red_tx_m_read_read                               : in  std_logic                     := 'X';             -- read
			red_tx_m_read_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			red_tx_m_read_readdatavalid                      : out std_logic;                                        -- readdatavalid
			ted_decryptor_read_master_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			ted_decryptor_read_master_waitrequest            : out std_logic;                                        -- waitrequest
			ted_decryptor_read_master_read                   : in  std_logic                     := 'X';             -- read
			ted_decryptor_read_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			ted_decryptor_write_master_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			ted_decryptor_write_master_waitrequest           : out std_logic;                                        -- waitrequest
			ted_decryptor_write_master_write                 : in  std_logic                     := 'X';             -- write
			ted_decryptor_write_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ted_encryptor_read_master_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			ted_encryptor_read_master_waitrequest            : out std_logic;                                        -- waitrequest
			ted_encryptor_read_master_read                   : in  std_logic                     := 'X';             -- read
			ted_encryptor_read_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			ted_encryptor_write_master_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			ted_encryptor_write_master_waitrequest           : out std_logic;                                        -- waitrequest
			ted_encryptor_write_master_write                 : in  std_logic                     := 'X';             -- write
			ted_encryptor_write_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			black_interface_control_port_address             : out std_logic_vector(7 downto 0);                     -- address
			black_interface_control_port_write               : out std_logic;                                        -- write
			black_interface_control_port_read                : out std_logic;                                        -- read
			black_interface_control_port_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			black_interface_control_port_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			black_interface_control_port_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			black_rx_csr_address                             : out std_logic_vector(3 downto 0);                     -- address
			black_rx_csr_write                               : out std_logic;                                        -- write
			black_rx_csr_read                                : out std_logic;                                        -- read
			black_rx_csr_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			black_rx_csr_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			black_rx_csr_chipselect                          : out std_logic;                                        -- chipselect
			black_to_red_memory_s1_address                   : out std_logic_vector(13 downto 0);                    -- address
			black_to_red_memory_s1_write                     : out std_logic;                                        -- write
			black_to_red_memory_s1_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			black_to_red_memory_s1_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			black_to_red_memory_s1_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			black_to_red_memory_s1_chipselect                : out std_logic;                                        -- chipselect
			black_to_red_memory_s1_clken                     : out std_logic;                                        -- clken
			black_tx_csr_address                             : out std_logic_vector(3 downto 0);                     -- address
			black_tx_csr_write                               : out std_logic;                                        -- write
			black_tx_csr_read                                : out std_logic;                                        -- read
			black_tx_csr_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			black_tx_csr_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			black_tx_csr_chipselect                          : out std_logic;                                        -- chipselect
			descriptor_mem_s1_address                        : out std_logic_vector(12 downto 0);                    -- address
			descriptor_mem_s1_write                          : out std_logic;                                        -- write
			descriptor_mem_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_mem_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_mem_s1_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_mem_s1_chipselect                     : out std_logic;                                        -- chipselect
			descriptor_mem_s1_clken                          : out std_logic;                                        -- clken
			heap_stack_s1_address                            : out std_logic_vector(12 downto 0);                    -- address
			heap_stack_s1_write                              : out std_logic;                                        -- write
			heap_stack_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			heap_stack_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			heap_stack_s1_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			heap_stack_s1_chipselect                         : out std_logic;                                        -- chipselect
			heap_stack_s1_clken                              : out std_logic;                                        -- clken
			hex_avalon_slave_0_write                         : out std_logic;                                        -- write
			hex_avalon_slave_0_read                          : out std_logic;                                        -- read
			hex_avalon_slave_0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			hex_avalon_slave_0_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			hex_avalon_slave_0_chipselect                    : out std_logic;                                        -- chipselect
			input_port_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			input_port_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			instruction_memory_s1_address                    : out std_logic_vector(15 downto 0);                    -- address
			instruction_memory_s1_write                      : out std_logic;                                        -- write
			instruction_memory_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			instruction_memory_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			instruction_memory_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			instruction_memory_s1_chipselect                 : out std_logic;                                        -- chipselect
			instruction_memory_s1_clken                      : out std_logic;                                        -- clken
			jtag_uart_avalon_jtag_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                 : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect           : out std_logic;                                        -- chipselect
			lcd_avalon_lcd_slave_address                     : out std_logic_vector(0 downto 0);                     -- address
			lcd_avalon_lcd_slave_write                       : out std_logic;                                        -- write
			lcd_avalon_lcd_slave_read                        : out std_logic;                                        -- read
			lcd_avalon_lcd_slave_readdata                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			lcd_avalon_lcd_slave_writedata                   : out std_logic_vector(7 downto 0);                     -- writedata
			lcd_avalon_lcd_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			lcd_avalon_lcd_slave_chipselect                  : out std_logic;                                        -- chipselect
			lcd_clk_pll_slave_address                        : out std_logic_vector(1 downto 0);                     -- address
			lcd_clk_pll_slave_write                          : out std_logic;                                        -- write
			lcd_clk_pll_slave_read                           : out std_logic;                                        -- read
			lcd_clk_pll_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lcd_clk_pll_slave_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_0_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_qsys_0_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_qsys_0_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_0_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			output_port_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			output_port_s1_write                             : out std_logic;                                        -- write
			output_port_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			output_port_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			output_port_s1_chipselect                        : out std_logic;                                        -- chipselect
			red_interface_control_port_address               : out std_logic_vector(7 downto 0);                     -- address
			red_interface_control_port_write                 : out std_logic;                                        -- write
			red_interface_control_port_read                  : out std_logic;                                        -- read
			red_interface_control_port_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			red_interface_control_port_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			red_interface_control_port_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			red_rx_csr_address                               : out std_logic_vector(3 downto 0);                     -- address
			red_rx_csr_write                                 : out std_logic;                                        -- write
			red_rx_csr_read                                  : out std_logic;                                        -- read
			red_rx_csr_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			red_rx_csr_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			red_rx_csr_chipselect                            : out std_logic;                                        -- chipselect
			red_to_black_memory_s1_address                   : out std_logic_vector(13 downto 0);                    -- address
			red_to_black_memory_s1_write                     : out std_logic;                                        -- write
			red_to_black_memory_s1_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			red_to_black_memory_s1_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			red_to_black_memory_s1_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			red_to_black_memory_s1_chipselect                : out std_logic;                                        -- chipselect
			red_to_black_memory_s1_clken                     : out std_logic;                                        -- clken
			red_tx_csr_address                               : out std_logic_vector(3 downto 0);                     -- address
			red_tx_csr_write                                 : out std_logic;                                        -- write
			red_tx_csr_read                                  : out std_logic;                                        -- read
			red_tx_csr_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			red_tx_csr_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			red_tx_csr_chipselect                            : out std_logic;                                        -- chipselect
			system_id_control_slave_address                  : out std_logic_vector(0 downto 0);                     -- address
			system_id_control_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			system_timer_s1_address                          : out std_logic_vector(3 downto 0);                     -- address
			system_timer_s1_write                            : out std_logic;                                        -- write
			system_timer_s1_readdata                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			system_timer_s1_writedata                        : out std_logic_vector(15 downto 0);                    -- writedata
			system_timer_s1_chipselect                       : out std_logic;                                        -- chipselect
			ted_decryptor_csr_address                        : out std_logic_vector(2 downto 0);                     -- address
			ted_decryptor_csr_write                          : out std_logic;                                        -- write
			ted_decryptor_csr_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ted_decryptor_csr_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			ted_encryptor_csr_address                        : out std_logic_vector(2 downto 0);                     -- address
			ted_encryptor_csr_write                          : out std_logic;                                        -- write
			ted_encryptor_csr_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ted_encryptor_csr_writedata                      : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component TEDv3_architecture_mm_interconnect_0;

	component TEDv3_architecture_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component TEDv3_architecture_irq_mapper;

	component TEDv3_architecture_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic                                         -- error
		);
	end component TEDv3_architecture_avalon_st_adapter;

	component TEDv3_architecture_avalon_st_adapter_002 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0)                      -- empty
		);
	end component TEDv3_architecture_avalon_st_adapter_002;

	component tedv3_architecture_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component tedv3_architecture_rst_controller;

	component tedv3_architecture_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component tedv3_architecture_rst_controller_001;

	signal lcd_clk_c0_clk                                                : std_logic;                     -- lcd_clk:c0 -> [lcd:clk, mm_interconnect_0:lcd_clk_c0_clk, rst_controller_001:clk]
	signal nios2_qsys_0_data_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_debugaccess                          : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	signal nios2_qsys_0_data_master_address                              : std_logic_vector(25 downto 0); -- nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	signal nios2_qsys_0_data_master_byteenable                           : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	signal nios2_qsys_0_data_master_read                                 : std_logic;                     -- nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	signal nios2_qsys_0_data_master_write                                : std_logic;                     -- nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	signal nios2_qsys_0_data_master_writedata                            : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	signal red_rx_descriptor_read_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_rx_descriptor_read_readdata -> red_rx:descriptor_read_readdata
	signal red_rx_descriptor_read_waitrequest                            : std_logic;                     -- mm_interconnect_0:red_rx_descriptor_read_waitrequest -> red_rx:descriptor_read_waitrequest
	signal red_rx_descriptor_read_address                                : std_logic_vector(31 downto 0); -- red_rx:descriptor_read_address -> mm_interconnect_0:red_rx_descriptor_read_address
	signal red_rx_descriptor_read_read                                   : std_logic;                     -- red_rx:descriptor_read_read -> mm_interconnect_0:red_rx_descriptor_read_read
	signal red_rx_descriptor_read_readdatavalid                          : std_logic;                     -- mm_interconnect_0:red_rx_descriptor_read_readdatavalid -> red_rx:descriptor_read_readdatavalid
	signal red_tx_descriptor_read_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_tx_descriptor_read_readdata -> red_tx:descriptor_read_readdata
	signal red_tx_descriptor_read_waitrequest                            : std_logic;                     -- mm_interconnect_0:red_tx_descriptor_read_waitrequest -> red_tx:descriptor_read_waitrequest
	signal red_tx_descriptor_read_address                                : std_logic_vector(31 downto 0); -- red_tx:descriptor_read_address -> mm_interconnect_0:red_tx_descriptor_read_address
	signal red_tx_descriptor_read_read                                   : std_logic;                     -- red_tx:descriptor_read_read -> mm_interconnect_0:red_tx_descriptor_read_read
	signal red_tx_descriptor_read_readdatavalid                          : std_logic;                     -- mm_interconnect_0:red_tx_descriptor_read_readdatavalid -> red_tx:descriptor_read_readdatavalid
	signal black_rx_descriptor_read_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:black_rx_descriptor_read_readdata -> black_rx:descriptor_read_readdata
	signal black_rx_descriptor_read_waitrequest                          : std_logic;                     -- mm_interconnect_0:black_rx_descriptor_read_waitrequest -> black_rx:descriptor_read_waitrequest
	signal black_rx_descriptor_read_address                              : std_logic_vector(31 downto 0); -- black_rx:descriptor_read_address -> mm_interconnect_0:black_rx_descriptor_read_address
	signal black_rx_descriptor_read_read                                 : std_logic;                     -- black_rx:descriptor_read_read -> mm_interconnect_0:black_rx_descriptor_read_read
	signal black_rx_descriptor_read_readdatavalid                        : std_logic;                     -- mm_interconnect_0:black_rx_descriptor_read_readdatavalid -> black_rx:descriptor_read_readdatavalid
	signal black_tx_descriptor_read_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:black_tx_descriptor_read_readdata -> black_tx:descriptor_read_readdata
	signal black_tx_descriptor_read_waitrequest                          : std_logic;                     -- mm_interconnect_0:black_tx_descriptor_read_waitrequest -> black_tx:descriptor_read_waitrequest
	signal black_tx_descriptor_read_address                              : std_logic_vector(31 downto 0); -- black_tx:descriptor_read_address -> mm_interconnect_0:black_tx_descriptor_read_address
	signal black_tx_descriptor_read_read                                 : std_logic;                     -- black_tx:descriptor_read_read -> mm_interconnect_0:black_tx_descriptor_read_read
	signal black_tx_descriptor_read_readdatavalid                        : std_logic;                     -- mm_interconnect_0:black_tx_descriptor_read_readdatavalid -> black_tx:descriptor_read_readdatavalid
	signal red_rx_descriptor_write_waitrequest                           : std_logic;                     -- mm_interconnect_0:red_rx_descriptor_write_waitrequest -> red_rx:descriptor_write_waitrequest
	signal red_rx_descriptor_write_address                               : std_logic_vector(31 downto 0); -- red_rx:descriptor_write_address -> mm_interconnect_0:red_rx_descriptor_write_address
	signal red_rx_descriptor_write_write                                 : std_logic;                     -- red_rx:descriptor_write_write -> mm_interconnect_0:red_rx_descriptor_write_write
	signal red_rx_descriptor_write_writedata                             : std_logic_vector(31 downto 0); -- red_rx:descriptor_write_writedata -> mm_interconnect_0:red_rx_descriptor_write_writedata
	signal red_tx_descriptor_write_waitrequest                           : std_logic;                     -- mm_interconnect_0:red_tx_descriptor_write_waitrequest -> red_tx:descriptor_write_waitrequest
	signal red_tx_descriptor_write_address                               : std_logic_vector(31 downto 0); -- red_tx:descriptor_write_address -> mm_interconnect_0:red_tx_descriptor_write_address
	signal red_tx_descriptor_write_write                                 : std_logic;                     -- red_tx:descriptor_write_write -> mm_interconnect_0:red_tx_descriptor_write_write
	signal red_tx_descriptor_write_writedata                             : std_logic_vector(31 downto 0); -- red_tx:descriptor_write_writedata -> mm_interconnect_0:red_tx_descriptor_write_writedata
	signal black_rx_descriptor_write_waitrequest                         : std_logic;                     -- mm_interconnect_0:black_rx_descriptor_write_waitrequest -> black_rx:descriptor_write_waitrequest
	signal black_rx_descriptor_write_address                             : std_logic_vector(31 downto 0); -- black_rx:descriptor_write_address -> mm_interconnect_0:black_rx_descriptor_write_address
	signal black_rx_descriptor_write_write                               : std_logic;                     -- black_rx:descriptor_write_write -> mm_interconnect_0:black_rx_descriptor_write_write
	signal black_rx_descriptor_write_writedata                           : std_logic_vector(31 downto 0); -- black_rx:descriptor_write_writedata -> mm_interconnect_0:black_rx_descriptor_write_writedata
	signal black_tx_descriptor_write_waitrequest                         : std_logic;                     -- mm_interconnect_0:black_tx_descriptor_write_waitrequest -> black_tx:descriptor_write_waitrequest
	signal black_tx_descriptor_write_address                             : std_logic_vector(31 downto 0); -- black_tx:descriptor_write_address -> mm_interconnect_0:black_tx_descriptor_write_address
	signal black_tx_descriptor_write_write                               : std_logic;                     -- black_tx:descriptor_write_write -> mm_interconnect_0:black_tx_descriptor_write_write
	signal black_tx_descriptor_write_writedata                           : std_logic_vector(31 downto 0); -- black_tx:descriptor_write_writedata -> mm_interconnect_0:black_tx_descriptor_write_writedata
	signal red_tx_m_read_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_tx_m_read_readdata -> red_tx:m_read_readdata
	signal red_tx_m_read_waitrequest                                     : std_logic;                     -- mm_interconnect_0:red_tx_m_read_waitrequest -> red_tx:m_read_waitrequest
	signal red_tx_m_read_address                                         : std_logic_vector(31 downto 0); -- red_tx:m_read_address -> mm_interconnect_0:red_tx_m_read_address
	signal red_tx_m_read_read                                            : std_logic;                     -- red_tx:m_read_read -> mm_interconnect_0:red_tx_m_read_read
	signal red_tx_m_read_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:red_tx_m_read_readdatavalid -> red_tx:m_read_readdatavalid
	signal black_rx_m_write_waitrequest                                  : std_logic;                     -- mm_interconnect_0:black_rx_m_write_waitrequest -> black_rx:m_write_waitrequest
	signal black_rx_m_write_address                                      : std_logic_vector(31 downto 0); -- black_rx:m_write_address -> mm_interconnect_0:black_rx_m_write_address
	signal black_rx_m_write_byteenable                                   : std_logic_vector(3 downto 0);  -- black_rx:m_write_byteenable -> mm_interconnect_0:black_rx_m_write_byteenable
	signal black_rx_m_write_write                                        : std_logic;                     -- black_rx:m_write_write -> mm_interconnect_0:black_rx_m_write_write
	signal black_rx_m_write_writedata                                    : std_logic_vector(31 downto 0); -- black_rx:m_write_writedata -> mm_interconnect_0:black_rx_m_write_writedata
	signal ted_decryptor_read_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:ted_decryptor_read_master_readdata -> ted_decryptor:avm_read_master_readdata
	signal ted_decryptor_read_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:ted_decryptor_read_master_waitrequest -> ted_decryptor:avm_read_master_waitrequest
	signal ted_decryptor_read_master_read                                : std_logic;                     -- ted_decryptor:avm_read_master_read -> mm_interconnect_0:ted_decryptor_read_master_read
	signal ted_decryptor_read_master_address                             : std_logic_vector(31 downto 0); -- ted_decryptor:avm_read_master_address -> mm_interconnect_0:ted_decryptor_read_master_address
	signal ted_decryptor_write_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:ted_decryptor_write_master_waitrequest -> ted_decryptor:avm_write_master_waitrequest
	signal ted_decryptor_write_master_address                            : std_logic_vector(31 downto 0); -- ted_decryptor:avm_write_master_address -> mm_interconnect_0:ted_decryptor_write_master_address
	signal ted_decryptor_write_master_write                              : std_logic;                     -- ted_decryptor:avm_write_master_write -> mm_interconnect_0:ted_decryptor_write_master_write
	signal ted_decryptor_write_master_writedata                          : std_logic_vector(31 downto 0); -- ted_decryptor:avm_write_master_writedata -> mm_interconnect_0:ted_decryptor_write_master_writedata
	signal black_tx_m_read_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:black_tx_m_read_readdata -> black_tx:m_read_readdata
	signal black_tx_m_read_waitrequest                                   : std_logic;                     -- mm_interconnect_0:black_tx_m_read_waitrequest -> black_tx:m_read_waitrequest
	signal black_tx_m_read_address                                       : std_logic_vector(31 downto 0); -- black_tx:m_read_address -> mm_interconnect_0:black_tx_m_read_address
	signal black_tx_m_read_read                                          : std_logic;                     -- black_tx:m_read_read -> mm_interconnect_0:black_tx_m_read_read
	signal black_tx_m_read_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:black_tx_m_read_readdatavalid -> black_tx:m_read_readdatavalid
	signal red_rx_m_write_waitrequest                                    : std_logic;                     -- mm_interconnect_0:red_rx_m_write_waitrequest -> red_rx:m_write_waitrequest
	signal red_rx_m_write_address                                        : std_logic_vector(31 downto 0); -- red_rx:m_write_address -> mm_interconnect_0:red_rx_m_write_address
	signal red_rx_m_write_byteenable                                     : std_logic_vector(3 downto 0);  -- red_rx:m_write_byteenable -> mm_interconnect_0:red_rx_m_write_byteenable
	signal red_rx_m_write_write                                          : std_logic;                     -- red_rx:m_write_write -> mm_interconnect_0:red_rx_m_write_write
	signal red_rx_m_write_writedata                                      : std_logic_vector(31 downto 0); -- red_rx:m_write_writedata -> mm_interconnect_0:red_rx_m_write_writedata
	signal ted_encryptor_read_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:ted_encryptor_read_master_readdata -> ted_encryptor:avm_read_master_readdata
	signal ted_encryptor_read_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:ted_encryptor_read_master_waitrequest -> ted_encryptor:avm_read_master_waitrequest
	signal ted_encryptor_read_master_read                                : std_logic;                     -- ted_encryptor:avm_read_master_read -> mm_interconnect_0:ted_encryptor_read_master_read
	signal ted_encryptor_read_master_address                             : std_logic_vector(31 downto 0); -- ted_encryptor:avm_read_master_address -> mm_interconnect_0:ted_encryptor_read_master_address
	signal ted_encryptor_write_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:ted_encryptor_write_master_waitrequest -> ted_encryptor:avm_write_master_waitrequest
	signal ted_encryptor_write_master_address                            : std_logic_vector(31 downto 0); -- ted_encryptor:avm_write_master_address -> mm_interconnect_0:ted_encryptor_write_master_address
	signal ted_encryptor_write_master_write                              : std_logic;                     -- ted_encryptor:avm_write_master_write -> mm_interconnect_0:ted_encryptor_write_master_write
	signal ted_encryptor_write_master_writedata                          : std_logic_vector(31 downto 0); -- ted_encryptor:avm_write_master_writedata -> mm_interconnect_0:ted_encryptor_write_master_writedata
	signal nios2_qsys_0_instruction_master_readdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_instruction_master_waitrequest                   : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                       : std_logic_vector(20 downto 0); -- nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	signal nios2_qsys_0_instruction_master_read                          : std_logic;                     -- nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_lcd_avalon_lcd_slave_chipselect             : std_logic;                     -- mm_interconnect_0:lcd_avalon_lcd_slave_chipselect -> lcd:chipselect
	signal mm_interconnect_0_lcd_avalon_lcd_slave_readdata               : std_logic_vector(7 downto 0);  -- lcd:readdata -> mm_interconnect_0:lcd_avalon_lcd_slave_readdata
	signal mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest            : std_logic;                     -- lcd:waitrequest -> mm_interconnect_0:lcd_avalon_lcd_slave_waitrequest
	signal mm_interconnect_0_lcd_avalon_lcd_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:lcd_avalon_lcd_slave_address -> lcd:address
	signal mm_interconnect_0_lcd_avalon_lcd_slave_read                   : std_logic;                     -- mm_interconnect_0:lcd_avalon_lcd_slave_read -> lcd:read
	signal mm_interconnect_0_lcd_avalon_lcd_slave_write                  : std_logic;                     -- mm_interconnect_0:lcd_avalon_lcd_slave_write -> lcd:write
	signal mm_interconnect_0_lcd_avalon_lcd_slave_writedata              : std_logic_vector(7 downto 0);  -- mm_interconnect_0:lcd_avalon_lcd_slave_writedata -> lcd:writedata
	signal mm_interconnect_0_hex_avalon_slave_0_chipselect               : std_logic;                     -- mm_interconnect_0:hex_avalon_slave_0_chipselect -> hex:chipselect
	signal mm_interconnect_0_hex_avalon_slave_0_readdata                 : std_logic_vector(31 downto 0); -- hex:readdata -> mm_interconnect_0:hex_avalon_slave_0_readdata
	signal mm_interconnect_0_hex_avalon_slave_0_read                     : std_logic;                     -- mm_interconnect_0:hex_avalon_slave_0_read -> hex:read
	signal mm_interconnect_0_hex_avalon_slave_0_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:hex_avalon_slave_0_byteenable -> hex:byteenable
	signal mm_interconnect_0_hex_avalon_slave_0_write                    : std_logic;                     -- mm_interconnect_0:hex_avalon_slave_0_write -> hex:write
	signal mm_interconnect_0_hex_avalon_slave_0_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_avalon_slave_0_writedata -> hex:writedata
	signal mm_interconnect_0_black_interface_control_port_readdata       : std_logic_vector(31 downto 0); -- black_interface:reg_data_out -> mm_interconnect_0:black_interface_control_port_readdata
	signal mm_interconnect_0_black_interface_control_port_waitrequest    : std_logic;                     -- black_interface:reg_busy -> mm_interconnect_0:black_interface_control_port_waitrequest
	signal mm_interconnect_0_black_interface_control_port_address        : std_logic_vector(7 downto 0);  -- mm_interconnect_0:black_interface_control_port_address -> black_interface:reg_addr
	signal mm_interconnect_0_black_interface_control_port_read           : std_logic;                     -- mm_interconnect_0:black_interface_control_port_read -> black_interface:reg_rd
	signal mm_interconnect_0_black_interface_control_port_write          : std_logic;                     -- mm_interconnect_0:black_interface_control_port_write -> black_interface:reg_wr
	signal mm_interconnect_0_black_interface_control_port_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:black_interface_control_port_writedata -> black_interface:reg_data_in
	signal mm_interconnect_0_red_interface_control_port_readdata         : std_logic_vector(31 downto 0); -- red_interface:reg_data_out -> mm_interconnect_0:red_interface_control_port_readdata
	signal mm_interconnect_0_red_interface_control_port_waitrequest      : std_logic;                     -- red_interface:reg_busy -> mm_interconnect_0:red_interface_control_port_waitrequest
	signal mm_interconnect_0_red_interface_control_port_address          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:red_interface_control_port_address -> red_interface:reg_addr
	signal mm_interconnect_0_red_interface_control_port_read             : std_logic;                     -- mm_interconnect_0:red_interface_control_port_read -> red_interface:reg_rd
	signal mm_interconnect_0_red_interface_control_port_write            : std_logic;                     -- mm_interconnect_0:red_interface_control_port_write -> red_interface:reg_wr
	signal mm_interconnect_0_red_interface_control_port_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_interface_control_port_writedata -> red_interface:reg_data_in
	signal mm_interconnect_0_system_id_control_slave_readdata            : std_logic_vector(31 downto 0); -- system_id:readdata -> mm_interconnect_0:system_id_control_slave_readdata
	signal mm_interconnect_0_system_id_control_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:system_id_control_slave_address -> system_id:address
	signal mm_interconnect_0_ted_encryptor_csr_readdata                  : std_logic_vector(31 downto 0); -- ted_encryptor:avs_csr_readdata -> mm_interconnect_0:ted_encryptor_csr_readdata
	signal mm_interconnect_0_ted_encryptor_csr_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ted_encryptor_csr_address -> ted_encryptor:avs_csr_address
	signal mm_interconnect_0_ted_encryptor_csr_write                     : std_logic;                     -- mm_interconnect_0:ted_encryptor_csr_write -> ted_encryptor:avs_csr_write
	signal mm_interconnect_0_ted_encryptor_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:ted_encryptor_csr_writedata -> ted_encryptor:avs_csr_writedata
	signal mm_interconnect_0_ted_decryptor_csr_readdata                  : std_logic_vector(31 downto 0); -- ted_decryptor:avs_csr_readdata -> mm_interconnect_0:ted_decryptor_csr_readdata
	signal mm_interconnect_0_ted_decryptor_csr_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ted_decryptor_csr_address -> ted_decryptor:avs_csr_address
	signal mm_interconnect_0_ted_decryptor_csr_write                     : std_logic;                     -- mm_interconnect_0:ted_decryptor_csr_write -> ted_decryptor:avs_csr_write
	signal mm_interconnect_0_ted_decryptor_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:ted_decryptor_csr_writedata -> ted_decryptor:avs_csr_writedata
	signal mm_interconnect_0_red_rx_csr_chipselect                       : std_logic;                     -- mm_interconnect_0:red_rx_csr_chipselect -> red_rx:csr_chipselect
	signal mm_interconnect_0_red_rx_csr_readdata                         : std_logic_vector(31 downto 0); -- red_rx:csr_readdata -> mm_interconnect_0:red_rx_csr_readdata
	signal mm_interconnect_0_red_rx_csr_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:red_rx_csr_address -> red_rx:csr_address
	signal mm_interconnect_0_red_rx_csr_read                             : std_logic;                     -- mm_interconnect_0:red_rx_csr_read -> red_rx:csr_read
	signal mm_interconnect_0_red_rx_csr_write                            : std_logic;                     -- mm_interconnect_0:red_rx_csr_write -> red_rx:csr_write
	signal mm_interconnect_0_red_rx_csr_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_rx_csr_writedata -> red_rx:csr_writedata
	signal mm_interconnect_0_red_tx_csr_chipselect                       : std_logic;                     -- mm_interconnect_0:red_tx_csr_chipselect -> red_tx:csr_chipselect
	signal mm_interconnect_0_red_tx_csr_readdata                         : std_logic_vector(31 downto 0); -- red_tx:csr_readdata -> mm_interconnect_0:red_tx_csr_readdata
	signal mm_interconnect_0_red_tx_csr_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:red_tx_csr_address -> red_tx:csr_address
	signal mm_interconnect_0_red_tx_csr_read                             : std_logic;                     -- mm_interconnect_0:red_tx_csr_read -> red_tx:csr_read
	signal mm_interconnect_0_red_tx_csr_write                            : std_logic;                     -- mm_interconnect_0:red_tx_csr_write -> red_tx:csr_write
	signal mm_interconnect_0_red_tx_csr_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_tx_csr_writedata -> red_tx:csr_writedata
	signal mm_interconnect_0_black_rx_csr_chipselect                     : std_logic;                     -- mm_interconnect_0:black_rx_csr_chipselect -> black_rx:csr_chipselect
	signal mm_interconnect_0_black_rx_csr_readdata                       : std_logic_vector(31 downto 0); -- black_rx:csr_readdata -> mm_interconnect_0:black_rx_csr_readdata
	signal mm_interconnect_0_black_rx_csr_address                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:black_rx_csr_address -> black_rx:csr_address
	signal mm_interconnect_0_black_rx_csr_read                           : std_logic;                     -- mm_interconnect_0:black_rx_csr_read -> black_rx:csr_read
	signal mm_interconnect_0_black_rx_csr_write                          : std_logic;                     -- mm_interconnect_0:black_rx_csr_write -> black_rx:csr_write
	signal mm_interconnect_0_black_rx_csr_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:black_rx_csr_writedata -> black_rx:csr_writedata
	signal mm_interconnect_0_black_tx_csr_chipselect                     : std_logic;                     -- mm_interconnect_0:black_tx_csr_chipselect -> black_tx:csr_chipselect
	signal mm_interconnect_0_black_tx_csr_readdata                       : std_logic_vector(31 downto 0); -- black_tx:csr_readdata -> mm_interconnect_0:black_tx_csr_readdata
	signal mm_interconnect_0_black_tx_csr_address                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:black_tx_csr_address -> black_tx:csr_address
	signal mm_interconnect_0_black_tx_csr_read                           : std_logic;                     -- mm_interconnect_0:black_tx_csr_read -> black_tx:csr_read
	signal mm_interconnect_0_black_tx_csr_write                          : std_logic;                     -- mm_interconnect_0:black_tx_csr_write -> black_tx:csr_write
	signal mm_interconnect_0_black_tx_csr_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:black_tx_csr_writedata -> black_tx:csr_writedata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata     : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest  : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess  : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address      : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read         : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write        : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal mm_interconnect_0_lcd_clk_pll_slave_readdata                  : std_logic_vector(31 downto 0); -- lcd_clk:readdata -> mm_interconnect_0:lcd_clk_pll_slave_readdata
	signal mm_interconnect_0_lcd_clk_pll_slave_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:lcd_clk_pll_slave_address -> lcd_clk:address
	signal mm_interconnect_0_lcd_clk_pll_slave_read                      : std_logic;                     -- mm_interconnect_0:lcd_clk_pll_slave_read -> lcd_clk:read
	signal mm_interconnect_0_lcd_clk_pll_slave_write                     : std_logic;                     -- mm_interconnect_0:lcd_clk_pll_slave_write -> lcd_clk:write
	signal mm_interconnect_0_lcd_clk_pll_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:lcd_clk_pll_slave_writedata -> lcd_clk:writedata
	signal mm_interconnect_0_output_port_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:output_port_s1_chipselect -> output_port:chipselect
	signal mm_interconnect_0_output_port_s1_readdata                     : std_logic_vector(31 downto 0); -- output_port:readdata -> mm_interconnect_0:output_port_s1_readdata
	signal mm_interconnect_0_output_port_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:output_port_s1_address -> output_port:address
	signal mm_interconnect_0_output_port_s1_write                        : std_logic;                     -- mm_interconnect_0:output_port_s1_write -> mm_interconnect_0_output_port_s1_write:in
	signal mm_interconnect_0_output_port_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:output_port_s1_writedata -> output_port:writedata
	signal mm_interconnect_0_input_port_s1_readdata                      : std_logic_vector(31 downto 0); -- input_port:readdata -> mm_interconnect_0:input_port_s1_readdata
	signal mm_interconnect_0_input_port_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:input_port_s1_address -> input_port:address
	signal mm_interconnect_0_instruction_memory_s1_chipselect            : std_logic;                     -- mm_interconnect_0:instruction_memory_s1_chipselect -> instruction_memory:chipselect
	signal mm_interconnect_0_instruction_memory_s1_readdata              : std_logic_vector(31 downto 0); -- instruction_memory:readdata -> mm_interconnect_0:instruction_memory_s1_readdata
	signal mm_interconnect_0_instruction_memory_s1_address               : std_logic_vector(15 downto 0); -- mm_interconnect_0:instruction_memory_s1_address -> instruction_memory:address
	signal mm_interconnect_0_instruction_memory_s1_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:instruction_memory_s1_byteenable -> instruction_memory:byteenable
	signal mm_interconnect_0_instruction_memory_s1_write                 : std_logic;                     -- mm_interconnect_0:instruction_memory_s1_write -> instruction_memory:write
	signal mm_interconnect_0_instruction_memory_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:instruction_memory_s1_writedata -> instruction_memory:writedata
	signal mm_interconnect_0_instruction_memory_s1_clken                 : std_logic;                     -- mm_interconnect_0:instruction_memory_s1_clken -> instruction_memory:clken
	signal mm_interconnect_0_heap_stack_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:heap_stack_s1_chipselect -> heap_stack:chipselect
	signal mm_interconnect_0_heap_stack_s1_readdata                      : std_logic_vector(31 downto 0); -- heap_stack:readdata -> mm_interconnect_0:heap_stack_s1_readdata
	signal mm_interconnect_0_heap_stack_s1_address                       : std_logic_vector(12 downto 0); -- mm_interconnect_0:heap_stack_s1_address -> heap_stack:address
	signal mm_interconnect_0_heap_stack_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:heap_stack_s1_byteenable -> heap_stack:byteenable
	signal mm_interconnect_0_heap_stack_s1_write                         : std_logic;                     -- mm_interconnect_0:heap_stack_s1_write -> heap_stack:write
	signal mm_interconnect_0_heap_stack_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:heap_stack_s1_writedata -> heap_stack:writedata
	signal mm_interconnect_0_heap_stack_s1_clken                         : std_logic;                     -- mm_interconnect_0:heap_stack_s1_clken -> heap_stack:clken
	signal mm_interconnect_0_system_timer_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:system_timer_s1_chipselect -> system_timer:chipselect
	signal mm_interconnect_0_system_timer_s1_readdata                    : std_logic_vector(15 downto 0); -- system_timer:readdata -> mm_interconnect_0:system_timer_s1_readdata
	signal mm_interconnect_0_system_timer_s1_address                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:system_timer_s1_address -> system_timer:address
	signal mm_interconnect_0_system_timer_s1_write                       : std_logic;                     -- mm_interconnect_0:system_timer_s1_write -> mm_interconnect_0_system_timer_s1_write:in
	signal mm_interconnect_0_system_timer_s1_writedata                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:system_timer_s1_writedata -> system_timer:writedata
	signal mm_interconnect_0_red_to_black_memory_s1_chipselect           : std_logic;                     -- mm_interconnect_0:red_to_black_memory_s1_chipselect -> red_to_black_memory:chipselect
	signal mm_interconnect_0_red_to_black_memory_s1_readdata             : std_logic_vector(31 downto 0); -- red_to_black_memory:readdata -> mm_interconnect_0:red_to_black_memory_s1_readdata
	signal mm_interconnect_0_red_to_black_memory_s1_address              : std_logic_vector(13 downto 0); -- mm_interconnect_0:red_to_black_memory_s1_address -> red_to_black_memory:address
	signal mm_interconnect_0_red_to_black_memory_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:red_to_black_memory_s1_byteenable -> red_to_black_memory:byteenable
	signal mm_interconnect_0_red_to_black_memory_s1_write                : std_logic;                     -- mm_interconnect_0:red_to_black_memory_s1_write -> red_to_black_memory:write
	signal mm_interconnect_0_red_to_black_memory_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_to_black_memory_s1_writedata -> red_to_black_memory:writedata
	signal mm_interconnect_0_red_to_black_memory_s1_clken                : std_logic;                     -- mm_interconnect_0:red_to_black_memory_s1_clken -> red_to_black_memory:clken
	signal mm_interconnect_0_black_to_red_memory_s1_chipselect           : std_logic;                     -- mm_interconnect_0:black_to_red_memory_s1_chipselect -> black_to_red_memory:chipselect
	signal mm_interconnect_0_black_to_red_memory_s1_readdata             : std_logic_vector(31 downto 0); -- black_to_red_memory:readdata -> mm_interconnect_0:black_to_red_memory_s1_readdata
	signal mm_interconnect_0_black_to_red_memory_s1_address              : std_logic_vector(13 downto 0); -- mm_interconnect_0:black_to_red_memory_s1_address -> black_to_red_memory:address
	signal mm_interconnect_0_black_to_red_memory_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:black_to_red_memory_s1_byteenable -> black_to_red_memory:byteenable
	signal mm_interconnect_0_black_to_red_memory_s1_write                : std_logic;                     -- mm_interconnect_0:black_to_red_memory_s1_write -> black_to_red_memory:write
	signal mm_interconnect_0_black_to_red_memory_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:black_to_red_memory_s1_writedata -> black_to_red_memory:writedata
	signal mm_interconnect_0_black_to_red_memory_s1_clken                : std_logic;                     -- mm_interconnect_0:black_to_red_memory_s1_clken -> black_to_red_memory:clken
	signal mm_interconnect_0_descriptor_mem_s1_chipselect                : std_logic;                     -- mm_interconnect_0:descriptor_mem_s1_chipselect -> descriptor_mem:chipselect
	signal mm_interconnect_0_descriptor_mem_s1_readdata                  : std_logic_vector(31 downto 0); -- descriptor_mem:readdata -> mm_interconnect_0:descriptor_mem_s1_readdata
	signal mm_interconnect_0_descriptor_mem_s1_address                   : std_logic_vector(12 downto 0); -- mm_interconnect_0:descriptor_mem_s1_address -> descriptor_mem:address
	signal mm_interconnect_0_descriptor_mem_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:descriptor_mem_s1_byteenable -> descriptor_mem:byteenable
	signal mm_interconnect_0_descriptor_mem_s1_write                     : std_logic;                     -- mm_interconnect_0:descriptor_mem_s1_write -> descriptor_mem:write
	signal mm_interconnect_0_descriptor_mem_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:descriptor_mem_s1_writedata -> descriptor_mem:writedata
	signal mm_interconnect_0_descriptor_mem_s1_clken                     : std_logic;                     -- mm_interconnect_0:descriptor_mem_s1_clken -> descriptor_mem:clken
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- red_rx:csr_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- red_tx:csr_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- black_rx:csr_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- black_tx:csr_irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                      : std_logic;                     -- system_timer:irq -> irq_mapper:receiver5_irq
	signal nios2_qsys_0_d_irq_irq                                        : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	signal black_tx_out_valid                                            : std_logic;                     -- black_tx:out_valid -> avalon_st_adapter:in_0_valid
	signal black_tx_out_data                                             : std_logic_vector(31 downto 0); -- black_tx:out_data -> avalon_st_adapter:in_0_data
	signal black_tx_out_ready                                            : std_logic;                     -- avalon_st_adapter:in_0_ready -> black_tx:out_ready
	signal black_tx_out_startofpacket                                    : std_logic;                     -- black_tx:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal black_tx_out_endofpacket                                      : std_logic;                     -- black_tx:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal black_tx_out_empty                                            : std_logic_vector(1 downto 0);  -- black_tx:out_empty -> avalon_st_adapter:in_0_empty
	signal avalon_st_adapter_out_0_valid                                 : std_logic;                     -- avalon_st_adapter:out_0_valid -> black_interface:ff_tx_wren
	signal avalon_st_adapter_out_0_data                                  : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> black_interface:ff_tx_data
	signal avalon_st_adapter_out_0_ready                                 : std_logic;                     -- black_interface:ff_tx_rdy -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                         : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> black_interface:ff_tx_sop
	signal avalon_st_adapter_out_0_endofpacket                           : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> black_interface:ff_tx_eop
	signal avalon_st_adapter_out_0_error                                 : std_logic;                     -- avalon_st_adapter:out_0_error -> black_interface:ff_tx_err
	signal avalon_st_adapter_out_0_empty                                 : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_empty -> black_interface:ff_tx_mod
	signal red_tx_out_valid                                              : std_logic;                     -- red_tx:out_valid -> avalon_st_adapter_001:in_0_valid
	signal red_tx_out_data                                               : std_logic_vector(31 downto 0); -- red_tx:out_data -> avalon_st_adapter_001:in_0_data
	signal red_tx_out_ready                                              : std_logic;                     -- avalon_st_adapter_001:in_0_ready -> red_tx:out_ready
	signal red_tx_out_startofpacket                                      : std_logic;                     -- red_tx:out_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	signal red_tx_out_endofpacket                                        : std_logic;                     -- red_tx:out_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	signal red_tx_out_empty                                              : std_logic_vector(1 downto 0);  -- red_tx:out_empty -> avalon_st_adapter_001:in_0_empty
	signal avalon_st_adapter_001_out_0_valid                             : std_logic;                     -- avalon_st_adapter_001:out_0_valid -> red_interface:ff_tx_wren
	signal avalon_st_adapter_001_out_0_data                              : std_logic_vector(31 downto 0); -- avalon_st_adapter_001:out_0_data -> red_interface:ff_tx_data
	signal avalon_st_adapter_001_out_0_ready                             : std_logic;                     -- red_interface:ff_tx_rdy -> avalon_st_adapter_001:out_0_ready
	signal avalon_st_adapter_001_out_0_startofpacket                     : std_logic;                     -- avalon_st_adapter_001:out_0_startofpacket -> red_interface:ff_tx_sop
	signal avalon_st_adapter_001_out_0_endofpacket                       : std_logic;                     -- avalon_st_adapter_001:out_0_endofpacket -> red_interface:ff_tx_eop
	signal avalon_st_adapter_001_out_0_error                             : std_logic;                     -- avalon_st_adapter_001:out_0_error -> red_interface:ff_tx_err
	signal avalon_st_adapter_001_out_0_empty                             : std_logic_vector(1 downto 0);  -- avalon_st_adapter_001:out_0_empty -> red_interface:ff_tx_mod
	signal black_interface_receive_valid                                 : std_logic;                     -- black_interface:ff_rx_dval -> avalon_st_adapter_002:in_0_valid
	signal black_interface_receive_data                                  : std_logic_vector(31 downto 0); -- black_interface:ff_rx_data -> avalon_st_adapter_002:in_0_data
	signal black_interface_receive_ready                                 : std_logic;                     -- avalon_st_adapter_002:in_0_ready -> black_interface:ff_rx_rdy
	signal black_interface_receive_startofpacket                         : std_logic;                     -- black_interface:ff_rx_sop -> avalon_st_adapter_002:in_0_startofpacket
	signal black_interface_receive_endofpacket                           : std_logic;                     -- black_interface:ff_rx_eop -> avalon_st_adapter_002:in_0_endofpacket
	signal black_interface_receive_error                                 : std_logic_vector(5 downto 0);  -- black_interface:rx_err -> avalon_st_adapter_002:in_0_error
	signal black_interface_receive_empty                                 : std_logic_vector(1 downto 0);  -- black_interface:ff_rx_mod -> avalon_st_adapter_002:in_0_empty
	signal avalon_st_adapter_002_out_0_valid                             : std_logic;                     -- avalon_st_adapter_002:out_0_valid -> black_rx:in_valid
	signal avalon_st_adapter_002_out_0_data                              : std_logic_vector(31 downto 0); -- avalon_st_adapter_002:out_0_data -> black_rx:in_data
	signal avalon_st_adapter_002_out_0_ready                             : std_logic;                     -- black_rx:in_ready -> avalon_st_adapter_002:out_0_ready
	signal avalon_st_adapter_002_out_0_startofpacket                     : std_logic;                     -- avalon_st_adapter_002:out_0_startofpacket -> black_rx:in_startofpacket
	signal avalon_st_adapter_002_out_0_endofpacket                       : std_logic;                     -- avalon_st_adapter_002:out_0_endofpacket -> black_rx:in_endofpacket
	signal avalon_st_adapter_002_out_0_empty                             : std_logic_vector(1 downto 0);  -- avalon_st_adapter_002:out_0_empty -> black_rx:in_empty
	signal red_interface_receive_valid                                   : std_logic;                     -- red_interface:ff_rx_dval -> avalon_st_adapter_003:in_0_valid
	signal red_interface_receive_data                                    : std_logic_vector(31 downto 0); -- red_interface:ff_rx_data -> avalon_st_adapter_003:in_0_data
	signal red_interface_receive_ready                                   : std_logic;                     -- avalon_st_adapter_003:in_0_ready -> red_interface:ff_rx_rdy
	signal red_interface_receive_startofpacket                           : std_logic;                     -- red_interface:ff_rx_sop -> avalon_st_adapter_003:in_0_startofpacket
	signal red_interface_receive_endofpacket                             : std_logic;                     -- red_interface:ff_rx_eop -> avalon_st_adapter_003:in_0_endofpacket
	signal red_interface_receive_error                                   : std_logic_vector(5 downto 0);  -- red_interface:rx_err -> avalon_st_adapter_003:in_0_error
	signal red_interface_receive_empty                                   : std_logic_vector(1 downto 0);  -- red_interface:ff_rx_mod -> avalon_st_adapter_003:in_0_empty
	signal avalon_st_adapter_003_out_0_valid                             : std_logic;                     -- avalon_st_adapter_003:out_0_valid -> red_rx:in_valid
	signal avalon_st_adapter_003_out_0_data                              : std_logic_vector(31 downto 0); -- avalon_st_adapter_003:out_0_data -> red_rx:in_data
	signal avalon_st_adapter_003_out_0_ready                             : std_logic;                     -- red_rx:in_ready -> avalon_st_adapter_003:out_0_ready
	signal avalon_st_adapter_003_out_0_startofpacket                     : std_logic;                     -- avalon_st_adapter_003:out_0_startofpacket -> red_rx:in_startofpacket
	signal avalon_st_adapter_003_out_0_endofpacket                       : std_logic;                     -- avalon_st_adapter_003:out_0_endofpacket -> red_rx:in_endofpacket
	signal avalon_st_adapter_003_out_0_empty                             : std_logic_vector(1 downto 0);  -- avalon_st_adapter_003:out_0_empty -> red_rx:in_empty
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, black_interface:reset, black_to_red_memory:reset, descriptor_mem:reset, heap_stack:reset, instruction_memory:reset, irq_mapper:reset, lcd_clk:reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, red_interface:reset, red_to_black_memory:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, ted_decryptor:csi_clock_reset, ted_encryptor:csi_clock_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [black_to_red_memory:reset_req, descriptor_mem:reset_req, heap_stack:reset_req, instruction_memory:reset_req, nios2_qsys_0:reset_req, red_to_black_memory:reset_req, rst_translator:reset_req_in]
	signal nios2_qsys_0_jtag_debug_module_reset_reset                    : std_logic;                     -- nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [lcd:reset, mm_interconnect_0:lcd_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_output_port_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_output_port_s1_write:inv -> output_port:write_n
	signal mm_interconnect_0_system_timer_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_0_system_timer_s1_write:inv -> system_timer:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [black_rx:system_reset_n, black_tx:system_reset_n, hex:resetn, input_port:reset_n, jtag_uart:rst_n, nios2_qsys_0:reset_n, output_port:reset_n, red_rx:system_reset_n, red_tx:system_reset_n, system_id:reset_n, system_timer:reset_n]

begin

	black_interface : component TEDv3_architecture_black_interface
		port map (
			clk           => clk_clk,                                                    -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                             --              reset_connection.reset
			reg_addr      => mm_interconnect_0_black_interface_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_0_black_interface_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_0_black_interface_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_0_black_interface_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_0_black_interface_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_0_black_interface_control_port_waitrequest, --                              .waitrequest
			tx_clk        => black_interface_pcs_mac_tx_clock_connection_clk,            --   pcs_mac_tx_clock_connection.clk
			rx_clk        => black_interface_pcs_mac_rx_clock_connection_clk,            --   pcs_mac_rx_clock_connection.clk
			set_10        => black_interface_mac_status_connection_set_10,               --         mac_status_connection.set_10
			set_1000      => black_interface_mac_status_connection_set_1000,             --                              .set_1000
			eth_mode      => black_interface_mac_status_connection_eth_mode,             --                              .eth_mode
			ena_10        => black_interface_mac_status_connection_ena_10,               --                              .ena_10
			rgmii_in      => black_interface_mac_rgmii_connection_rgmii_in,              --          mac_rgmii_connection.rgmii_in
			rgmii_out     => black_interface_mac_rgmii_connection_rgmii_out,             --                              .rgmii_out
			rx_control    => black_interface_mac_rgmii_connection_rx_control,            --                              .rx_control
			tx_control    => black_interface_mac_rgmii_connection_tx_control,            --                              .tx_control
			ff_rx_clk     => clk_clk,                                                    --      receive_clock_connection.clk
			ff_tx_clk     => clk_clk,                                                    --     transmit_clock_connection.clk
			ff_rx_data    => black_interface_receive_data,                               --                       receive.data
			ff_rx_eop     => black_interface_receive_endofpacket,                        --                              .endofpacket
			rx_err        => black_interface_receive_error,                              --                              .error
			ff_rx_mod     => black_interface_receive_empty,                              --                              .empty
			ff_rx_rdy     => black_interface_receive_ready,                              --                              .ready
			ff_rx_sop     => black_interface_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => black_interface_receive_valid,                              --                              .valid
			ff_tx_data    => avalon_st_adapter_out_0_data,                               --                      transmit.data
			ff_tx_eop     => avalon_st_adapter_out_0_endofpacket,                        --                              .endofpacket
			ff_tx_err     => avalon_st_adapter_out_0_error,                              --                              .error
			ff_tx_mod     => avalon_st_adapter_out_0_empty,                              --                              .empty
			ff_tx_rdy     => avalon_st_adapter_out_0_ready,                              --                              .ready
			ff_tx_sop     => avalon_st_adapter_out_0_startofpacket,                      --                              .startofpacket
			ff_tx_wren    => avalon_st_adapter_out_0_valid,                              --                              .valid
			mdc           => black_interface_mac_mdio_connection_mdc,                    --           mac_mdio_connection.mdc
			mdio_in       => black_interface_mac_mdio_connection_mdio_in,                --                              .mdio_in
			mdio_out      => black_interface_mac_mdio_connection_mdio_out,               --                              .mdio_out
			mdio_oen      => black_interface_mac_mdio_connection_mdio_oen,               --                              .mdio_oen
			xon_gen       => black_interface_mac_misc_connection_xon_gen,                --           mac_misc_connection.xon_gen
			xoff_gen      => black_interface_mac_misc_connection_xoff_gen,               --                              .xoff_gen
			ff_tx_crc_fwd => black_interface_mac_misc_connection_ff_tx_crc_fwd,          --                              .ff_tx_crc_fwd
			ff_tx_septy   => black_interface_mac_misc_connection_ff_tx_septy,            --                              .ff_tx_septy
			tx_ff_uflow   => black_interface_mac_misc_connection_tx_ff_uflow,            --                              .tx_ff_uflow
			ff_tx_a_full  => black_interface_mac_misc_connection_ff_tx_a_full,           --                              .ff_tx_a_full
			ff_tx_a_empty => black_interface_mac_misc_connection_ff_tx_a_empty,          --                              .ff_tx_a_empty
			rx_err_stat   => black_interface_mac_misc_connection_rx_err_stat,            --                              .rx_err_stat
			rx_frm_type   => black_interface_mac_misc_connection_rx_frm_type,            --                              .rx_frm_type
			ff_rx_dsav    => black_interface_mac_misc_connection_ff_rx_dsav,             --                              .ff_rx_dsav
			ff_rx_a_full  => black_interface_mac_misc_connection_ff_rx_a_full,           --                              .ff_rx_a_full
			ff_rx_a_empty => black_interface_mac_misc_connection_ff_rx_a_empty           --                              .ff_rx_a_empty
		);

	black_rx : component TEDv3_architecture_black_rx
		port map (
			clk                           => clk_clk,                                   --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_black_rx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_black_rx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_black_rx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_black_rx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_black_rx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_black_rx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => black_rx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => black_rx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => black_rx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => black_rx_descriptor_read_address,          --                 .address
			descriptor_read_read          => black_rx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => black_rx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => black_rx_descriptor_write_address,         --                 .address
			descriptor_write_write        => black_rx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => black_rx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver2_irq,                  --          csr_irq.irq
			in_startofpacket              => avalon_st_adapter_002_out_0_startofpacket, --               in.startofpacket
			in_endofpacket                => avalon_st_adapter_002_out_0_endofpacket,   --                 .endofpacket
			in_data                       => avalon_st_adapter_002_out_0_data,          --                 .data
			in_valid                      => avalon_st_adapter_002_out_0_valid,         --                 .valid
			in_ready                      => avalon_st_adapter_002_out_0_ready,         --                 .ready
			in_empty                      => avalon_st_adapter_002_out_0_empty,         --                 .empty
			m_write_waitrequest           => black_rx_m_write_waitrequest,              --          m_write.waitrequest
			m_write_address               => black_rx_m_write_address,                  --                 .address
			m_write_write                 => black_rx_m_write_write,                    --                 .write
			m_write_writedata             => black_rx_m_write_writedata,                --                 .writedata
			m_write_byteenable            => black_rx_m_write_byteenable                --                 .byteenable
		);

	black_to_red_memory : component TEDv3_architecture_black_to_red_memory
		port map (
			clk        => clk_clk,                                             --   clk1.clk
			address    => mm_interconnect_0_black_to_red_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_black_to_red_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_black_to_red_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_black_to_red_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_black_to_red_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_black_to_red_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_black_to_red_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                   --       .reset_req
		);

	black_tx : component TEDv3_architecture_black_tx
		port map (
			clk                           => clk_clk,                                   --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_black_tx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_black_tx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_black_tx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_black_tx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_black_tx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_black_tx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => black_tx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => black_tx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => black_tx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => black_tx_descriptor_read_address,          --                 .address
			descriptor_read_read          => black_tx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => black_tx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => black_tx_descriptor_write_address,         --                 .address
			descriptor_write_write        => black_tx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => black_tx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver3_irq,                  --          csr_irq.irq
			m_read_readdata               => black_tx_m_read_readdata,                  --           m_read.readdata
			m_read_readdatavalid          => black_tx_m_read_readdatavalid,             --                 .readdatavalid
			m_read_waitrequest            => black_tx_m_read_waitrequest,               --                 .waitrequest
			m_read_address                => black_tx_m_read_address,                   --                 .address
			m_read_read                   => black_tx_m_read_read,                      --                 .read
			out_data                      => black_tx_out_data,                         --              out.data
			out_valid                     => black_tx_out_valid,                        --                 .valid
			out_ready                     => black_tx_out_ready,                        --                 .ready
			out_endofpacket               => black_tx_out_endofpacket,                  --                 .endofpacket
			out_startofpacket             => black_tx_out_startofpacket,                --                 .startofpacket
			out_empty                     => black_tx_out_empty                         --                 .empty
		);

	descriptor_mem : component TEDv3_architecture_descriptor_mem
		port map (
			clk        => clk_clk,                                        --   clk1.clk
			address    => mm_interconnect_0_descriptor_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_descriptor_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_descriptor_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_descriptor_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_descriptor_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_descriptor_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_descriptor_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req              --       .reset_req
		);

	heap_stack : component TEDv3_architecture_heap_stack
		port map (
			clk        => clk_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_heap_stack_s1_address,    --     s1.address
			clken      => mm_interconnect_0_heap_stack_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_heap_stack_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_heap_stack_s1_write,      --       .write
			readdata   => mm_interconnect_0_heap_stack_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_heap_stack_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_heap_stack_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req          --       .reset_req
		);

	hex : component reg32_avalon_interface
		port map (
			read       => mm_interconnect_0_hex_avalon_slave_0_read,       -- avalon_slave_0.read
			write      => mm_interconnect_0_hex_avalon_slave_0_write,      --               .write
			chipselect => mm_interconnect_0_hex_avalon_slave_0_chipselect, --               .chipselect
			writedata  => mm_interconnect_0_hex_avalon_slave_0_writedata,  --               .writedata
			byteenable => mm_interconnect_0_hex_avalon_slave_0_byteenable, --               .byteenable
			readdata   => mm_interconnect_0_hex_avalon_slave_0_readdata,   --               .readdata
			clock      => clk_clk,                                         --     clock_sink.clk
			resetn     => rst_controller_reset_out_reset_ports_inv,        --     reset_sink.reset_n
			Q_export   => hex_conduit_hex_conduit                          --    conduit_end.hex_conduit
		);

	input_port : component TEDv3_architecture_input_port
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_input_port_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_input_port_s1_readdata, --                    .readdata
			in_port  => input_port_external_connection_export     -- external_connection.export
		);

	instruction_memory : component TEDv3_architecture_instruction_memory
		port map (
			clk        => clk_clk,                                            --   clk1.clk
			address    => mm_interconnect_0_instruction_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_instruction_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_instruction_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_instruction_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_instruction_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_instruction_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_instruction_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                     -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                  --       .reset_req
		);

	jtag_uart : component TEDv3_architecture_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver4_irq                                       --               irq.irq
		);

	lcd : component TEDv3_architecture_lcd
		port map (
			clk         => lcd_clk_c0_clk,                                     --                clk.clk
			reset       => rst_controller_001_reset_out_reset,                 --              reset.reset
			address     => mm_interconnect_0_lcd_avalon_lcd_slave_address(0),  --   avalon_lcd_slave.address
			chipselect  => mm_interconnect_0_lcd_avalon_lcd_slave_chipselect,  --                   .chipselect
			read        => mm_interconnect_0_lcd_avalon_lcd_slave_read,        --                   .read
			write       => mm_interconnect_0_lcd_avalon_lcd_slave_write,       --                   .write
			writedata   => mm_interconnect_0_lcd_avalon_lcd_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_lcd_avalon_lcd_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest, --                   .waitrequest
			LCD_DATA    => lcd_external_interface_DATA,                        -- external_interface.export
			LCD_ON      => lcd_external_interface_ON,                          --                   .export
			LCD_BLON    => lcd_external_interface_BLON,                        --                   .export
			LCD_EN      => lcd_external_interface_EN,                          --                   .export
			LCD_RS      => lcd_external_interface_RS,                          --                   .export
			LCD_RW      => lcd_external_interface_RW                           --                   .export
		);

	lcd_clk : component TEDv3_architecture_lcd_clk
		port map (
			clk       => clk_clk,                                       --       inclk_interface.clk
			reset     => rst_controller_reset_out_reset,                -- inclk_interface_reset.reset
			read      => mm_interconnect_0_lcd_clk_pll_slave_read,      --             pll_slave.read
			write     => mm_interconnect_0_lcd_clk_pll_slave_write,     --                      .write
			address   => mm_interconnect_0_lcd_clk_pll_slave_address,   --                      .address
			readdata  => mm_interconnect_0_lcd_clk_pll_slave_readdata,  --                      .readdata
			writedata => mm_interconnect_0_lcd_clk_pll_slave_writedata, --                      .writedata
			c0        => lcd_clk_c0_clk,                                --                    c0.clk
			areset    => lcd_clk_areset_conduit_export,                 --        areset_conduit.export
			locked    => lcd_clk_locked_conduit_export,                 --        locked_conduit.export
			phasedone => lcd_clk_phasedone_conduit_export               --     phasedone_conduit.export
		);

	nios2_qsys_0 : component TEDv3_architecture_nios2_qsys_0
		port map (
			clk                                   => clk_clk,                                                      --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                     --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                           --                          .reset_req
			d_address                             => nios2_qsys_0_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_0_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                          -- custom_instruction_master.readra
		);

	output_port : component TEDv3_architecture_output_port
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_output_port_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_output_port_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_output_port_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_output_port_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_output_port_s1_readdata,        --                    .readdata
			out_port   => output_port_external_connection_export            -- external_connection.export
		);

	red_interface : component TEDv3_architecture_black_interface
		port map (
			clk           => clk_clk,                                                  -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                           --              reset_connection.reset
			reg_addr      => mm_interconnect_0_red_interface_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_0_red_interface_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_0_red_interface_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_0_red_interface_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_0_red_interface_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_0_red_interface_control_port_waitrequest, --                              .waitrequest
			tx_clk        => red_interface_pcs_mac_tx_clock_connection_clk,            --   pcs_mac_tx_clock_connection.clk
			rx_clk        => red_interface_pcs_mac_rx_clock_connection_clk,            --   pcs_mac_rx_clock_connection.clk
			set_10        => red_interface_mac_status_connection_set_10,               --         mac_status_connection.set_10
			set_1000      => red_interface_mac_status_connection_set_1000,             --                              .set_1000
			eth_mode      => red_interface_mac_status_connection_eth_mode,             --                              .eth_mode
			ena_10        => red_interface_mac_status_connection_ena_10,               --                              .ena_10
			rgmii_in      => red_interface_mac_rgmii_connection_rgmii_in,              --          mac_rgmii_connection.rgmii_in
			rgmii_out     => red_interface_mac_rgmii_connection_rgmii_out,             --                              .rgmii_out
			rx_control    => red_interface_mac_rgmii_connection_rx_control,            --                              .rx_control
			tx_control    => red_interface_mac_rgmii_connection_tx_control,            --                              .tx_control
			ff_rx_clk     => clk_clk,                                                  --      receive_clock_connection.clk
			ff_tx_clk     => clk_clk,                                                  --     transmit_clock_connection.clk
			ff_rx_data    => red_interface_receive_data,                               --                       receive.data
			ff_rx_eop     => red_interface_receive_endofpacket,                        --                              .endofpacket
			rx_err        => red_interface_receive_error,                              --                              .error
			ff_rx_mod     => red_interface_receive_empty,                              --                              .empty
			ff_rx_rdy     => red_interface_receive_ready,                              --                              .ready
			ff_rx_sop     => red_interface_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => red_interface_receive_valid,                              --                              .valid
			ff_tx_data    => avalon_st_adapter_001_out_0_data,                         --                      transmit.data
			ff_tx_eop     => avalon_st_adapter_001_out_0_endofpacket,                  --                              .endofpacket
			ff_tx_err     => avalon_st_adapter_001_out_0_error,                        --                              .error
			ff_tx_mod     => avalon_st_adapter_001_out_0_empty,                        --                              .empty
			ff_tx_rdy     => avalon_st_adapter_001_out_0_ready,                        --                              .ready
			ff_tx_sop     => avalon_st_adapter_001_out_0_startofpacket,                --                              .startofpacket
			ff_tx_wren    => avalon_st_adapter_001_out_0_valid,                        --                              .valid
			mdc           => red_interface_mac_mdio_connection_mdc,                    --           mac_mdio_connection.mdc
			mdio_in       => red_interface_mac_mdio_connection_mdio_in,                --                              .mdio_in
			mdio_out      => red_interface_mac_mdio_connection_mdio_out,               --                              .mdio_out
			mdio_oen      => red_interface_mac_mdio_connection_mdio_oen,               --                              .mdio_oen
			xon_gen       => red_interface_mac_misc_connection_xon_gen,                --           mac_misc_connection.xon_gen
			xoff_gen      => red_interface_mac_misc_connection_xoff_gen,               --                              .xoff_gen
			ff_tx_crc_fwd => red_interface_mac_misc_connection_ff_tx_crc_fwd,          --                              .ff_tx_crc_fwd
			ff_tx_septy   => red_interface_mac_misc_connection_ff_tx_septy,            --                              .ff_tx_septy
			tx_ff_uflow   => red_interface_mac_misc_connection_tx_ff_uflow,            --                              .tx_ff_uflow
			ff_tx_a_full  => red_interface_mac_misc_connection_ff_tx_a_full,           --                              .ff_tx_a_full
			ff_tx_a_empty => red_interface_mac_misc_connection_ff_tx_a_empty,          --                              .ff_tx_a_empty
			rx_err_stat   => red_interface_mac_misc_connection_rx_err_stat,            --                              .rx_err_stat
			rx_frm_type   => red_interface_mac_misc_connection_rx_frm_type,            --                              .rx_frm_type
			ff_rx_dsav    => red_interface_mac_misc_connection_ff_rx_dsav,             --                              .ff_rx_dsav
			ff_rx_a_full  => red_interface_mac_misc_connection_ff_rx_a_full,           --                              .ff_rx_a_full
			ff_rx_a_empty => red_interface_mac_misc_connection_ff_rx_a_empty           --                              .ff_rx_a_empty
		);

	red_rx : component TEDv3_architecture_black_rx
		port map (
			clk                           => clk_clk,                                   --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_red_rx_csr_chipselect,   --              csr.chipselect
			csr_address                   => mm_interconnect_0_red_rx_csr_address,      --                 .address
			csr_read                      => mm_interconnect_0_red_rx_csr_read,         --                 .read
			csr_write                     => mm_interconnect_0_red_rx_csr_write,        --                 .write
			csr_writedata                 => mm_interconnect_0_red_rx_csr_writedata,    --                 .writedata
			csr_readdata                  => mm_interconnect_0_red_rx_csr_readdata,     --                 .readdata
			descriptor_read_readdata      => red_rx_descriptor_read_readdata,           --  descriptor_read.readdata
			descriptor_read_readdatavalid => red_rx_descriptor_read_readdatavalid,      --                 .readdatavalid
			descriptor_read_waitrequest   => red_rx_descriptor_read_waitrequest,        --                 .waitrequest
			descriptor_read_address       => red_rx_descriptor_read_address,            --                 .address
			descriptor_read_read          => red_rx_descriptor_read_read,               --                 .read
			descriptor_write_waitrequest  => red_rx_descriptor_write_waitrequest,       -- descriptor_write.waitrequest
			descriptor_write_address      => red_rx_descriptor_write_address,           --                 .address
			descriptor_write_write        => red_rx_descriptor_write_write,             --                 .write
			descriptor_write_writedata    => red_rx_descriptor_write_writedata,         --                 .writedata
			csr_irq                       => irq_mapper_receiver0_irq,                  --          csr_irq.irq
			in_startofpacket              => avalon_st_adapter_003_out_0_startofpacket, --               in.startofpacket
			in_endofpacket                => avalon_st_adapter_003_out_0_endofpacket,   --                 .endofpacket
			in_data                       => avalon_st_adapter_003_out_0_data,          --                 .data
			in_valid                      => avalon_st_adapter_003_out_0_valid,         --                 .valid
			in_ready                      => avalon_st_adapter_003_out_0_ready,         --                 .ready
			in_empty                      => avalon_st_adapter_003_out_0_empty,         --                 .empty
			m_write_waitrequest           => red_rx_m_write_waitrequest,                --          m_write.waitrequest
			m_write_address               => red_rx_m_write_address,                    --                 .address
			m_write_write                 => red_rx_m_write_write,                      --                 .write
			m_write_writedata             => red_rx_m_write_writedata,                  --                 .writedata
			m_write_byteenable            => red_rx_m_write_byteenable                  --                 .byteenable
		);

	red_to_black_memory : component TEDv3_architecture_red_to_black_memory
		port map (
			clk        => clk_clk,                                             --   clk1.clk
			address    => mm_interconnect_0_red_to_black_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_red_to_black_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_red_to_black_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_red_to_black_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_red_to_black_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_red_to_black_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_red_to_black_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                   --       .reset_req
		);

	red_tx : component TEDv3_architecture_black_tx
		port map (
			clk                           => clk_clk,                                  --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv, --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_red_tx_csr_chipselect,  --              csr.chipselect
			csr_address                   => mm_interconnect_0_red_tx_csr_address,     --                 .address
			csr_read                      => mm_interconnect_0_red_tx_csr_read,        --                 .read
			csr_write                     => mm_interconnect_0_red_tx_csr_write,       --                 .write
			csr_writedata                 => mm_interconnect_0_red_tx_csr_writedata,   --                 .writedata
			csr_readdata                  => mm_interconnect_0_red_tx_csr_readdata,    --                 .readdata
			descriptor_read_readdata      => red_tx_descriptor_read_readdata,          --  descriptor_read.readdata
			descriptor_read_readdatavalid => red_tx_descriptor_read_readdatavalid,     --                 .readdatavalid
			descriptor_read_waitrequest   => red_tx_descriptor_read_waitrequest,       --                 .waitrequest
			descriptor_read_address       => red_tx_descriptor_read_address,           --                 .address
			descriptor_read_read          => red_tx_descriptor_read_read,              --                 .read
			descriptor_write_waitrequest  => red_tx_descriptor_write_waitrequest,      -- descriptor_write.waitrequest
			descriptor_write_address      => red_tx_descriptor_write_address,          --                 .address
			descriptor_write_write        => red_tx_descriptor_write_write,            --                 .write
			descriptor_write_writedata    => red_tx_descriptor_write_writedata,        --                 .writedata
			csr_irq                       => irq_mapper_receiver1_irq,                 --          csr_irq.irq
			m_read_readdata               => red_tx_m_read_readdata,                   --           m_read.readdata
			m_read_readdatavalid          => red_tx_m_read_readdatavalid,              --                 .readdatavalid
			m_read_waitrequest            => red_tx_m_read_waitrequest,                --                 .waitrequest
			m_read_address                => red_tx_m_read_address,                    --                 .address
			m_read_read                   => red_tx_m_read_read,                       --                 .read
			out_data                      => red_tx_out_data,                          --              out.data
			out_valid                     => red_tx_out_valid,                         --                 .valid
			out_ready                     => red_tx_out_ready,                         --                 .ready
			out_endofpacket               => red_tx_out_endofpacket,                   --                 .endofpacket
			out_startofpacket             => red_tx_out_startofpacket,                 --                 .startofpacket
			out_empty                     => red_tx_out_empty                          --                 .empty
		);

	system_id : component TEDv3_architecture_system_id
		port map (
			clock    => clk_clk,                                              --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,             --         reset.reset_n
			readdata => mm_interconnect_0_system_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_system_id_control_slave_address(0)  --              .address
		);

	system_timer : component TEDv3_architecture_system_timer
		port map (
			clk        => clk_clk,                                           --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          -- reset.reset_n
			address    => mm_interconnect_0_system_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_system_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_system_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_system_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_system_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                           --   irq.irq
		);

	ted_decryptor : component ted_crypto
		port map (
			csi_clock_clk                => clk_clk,                                       --        clock.clk
			csi_clock_reset              => rst_controller_reset_out_reset,                --  clock_reset.reset
			avm_read_master_read         => ted_decryptor_read_master_read,                --  read_master.read
			avm_read_master_address      => ted_decryptor_read_master_address,             --             .address
			avm_read_master_readdata     => ted_decryptor_read_master_readdata,            --             .readdata
			avm_read_master_waitrequest  => ted_decryptor_read_master_waitrequest,         --             .waitrequest
			avm_write_master_write       => ted_decryptor_write_master_write,              -- write_master.write
			avm_write_master_address     => ted_decryptor_write_master_address,            --             .address
			avm_write_master_writedata   => ted_decryptor_write_master_writedata,          --             .writedata
			avm_write_master_waitrequest => ted_decryptor_write_master_waitrequest,        --             .waitrequest
			avs_csr_address              => mm_interconnect_0_ted_decryptor_csr_address,   --          csr.address
			avs_csr_readdata             => mm_interconnect_0_ted_decryptor_csr_readdata,  --             .readdata
			avs_csr_write                => mm_interconnect_0_ted_decryptor_csr_write,     --             .write
			avs_csr_writedata            => mm_interconnect_0_ted_decryptor_csr_writedata  --             .writedata
		);

	ted_encryptor : component ted_crypto
		port map (
			csi_clock_clk                => clk_clk,                                       --        clock.clk
			csi_clock_reset              => rst_controller_reset_out_reset,                --  clock_reset.reset
			avm_read_master_read         => ted_encryptor_read_master_read,                --  read_master.read
			avm_read_master_address      => ted_encryptor_read_master_address,             --             .address
			avm_read_master_readdata     => ted_encryptor_read_master_readdata,            --             .readdata
			avm_read_master_waitrequest  => ted_encryptor_read_master_waitrequest,         --             .waitrequest
			avm_write_master_write       => ted_encryptor_write_master_write,              -- write_master.write
			avm_write_master_address     => ted_encryptor_write_master_address,            --             .address
			avm_write_master_writedata   => ted_encryptor_write_master_writedata,          --             .writedata
			avm_write_master_waitrequest => ted_encryptor_write_master_waitrequest,        --             .waitrequest
			avs_csr_address              => mm_interconnect_0_ted_encryptor_csr_address,   --          csr.address
			avs_csr_readdata             => mm_interconnect_0_ted_encryptor_csr_readdata,  --             .readdata
			avs_csr_write                => mm_interconnect_0_ted_encryptor_csr_write,     --             .write
			avs_csr_writedata            => mm_interconnect_0_ted_encryptor_csr_writedata  --             .writedata
		);

	mm_interconnect_0 : component TEDv3_architecture_mm_interconnect_0
		port map (
			lcd_clk_c0_clk                                   => lcd_clk_c0_clk,                                               --                                 lcd_clk_c0.clk
			sys_clk_clk_clk                                  => clk_clk,                                                      --                                sys_clk_clk.clk
			lcd_reset_reset_bridge_in_reset_reset            => rst_controller_001_reset_out_reset,                           --            lcd_reset_reset_bridge_in_reset.reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                               -- nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
			black_rx_descriptor_read_address                 => black_rx_descriptor_read_address,                             --                   black_rx_descriptor_read.address
			black_rx_descriptor_read_waitrequest             => black_rx_descriptor_read_waitrequest,                         --                                           .waitrequest
			black_rx_descriptor_read_read                    => black_rx_descriptor_read_read,                                --                                           .read
			black_rx_descriptor_read_readdata                => black_rx_descriptor_read_readdata,                            --                                           .readdata
			black_rx_descriptor_read_readdatavalid           => black_rx_descriptor_read_readdatavalid,                       --                                           .readdatavalid
			black_rx_descriptor_write_address                => black_rx_descriptor_write_address,                            --                  black_rx_descriptor_write.address
			black_rx_descriptor_write_waitrequest            => black_rx_descriptor_write_waitrequest,                        --                                           .waitrequest
			black_rx_descriptor_write_write                  => black_rx_descriptor_write_write,                              --                                           .write
			black_rx_descriptor_write_writedata              => black_rx_descriptor_write_writedata,                          --                                           .writedata
			black_rx_m_write_address                         => black_rx_m_write_address,                                     --                           black_rx_m_write.address
			black_rx_m_write_waitrequest                     => black_rx_m_write_waitrequest,                                 --                                           .waitrequest
			black_rx_m_write_byteenable                      => black_rx_m_write_byteenable,                                  --                                           .byteenable
			black_rx_m_write_write                           => black_rx_m_write_write,                                       --                                           .write
			black_rx_m_write_writedata                       => black_rx_m_write_writedata,                                   --                                           .writedata
			black_tx_descriptor_read_address                 => black_tx_descriptor_read_address,                             --                   black_tx_descriptor_read.address
			black_tx_descriptor_read_waitrequest             => black_tx_descriptor_read_waitrequest,                         --                                           .waitrequest
			black_tx_descriptor_read_read                    => black_tx_descriptor_read_read,                                --                                           .read
			black_tx_descriptor_read_readdata                => black_tx_descriptor_read_readdata,                            --                                           .readdata
			black_tx_descriptor_read_readdatavalid           => black_tx_descriptor_read_readdatavalid,                       --                                           .readdatavalid
			black_tx_descriptor_write_address                => black_tx_descriptor_write_address,                            --                  black_tx_descriptor_write.address
			black_tx_descriptor_write_waitrequest            => black_tx_descriptor_write_waitrequest,                        --                                           .waitrequest
			black_tx_descriptor_write_write                  => black_tx_descriptor_write_write,                              --                                           .write
			black_tx_descriptor_write_writedata              => black_tx_descriptor_write_writedata,                          --                                           .writedata
			black_tx_m_read_address                          => black_tx_m_read_address,                                      --                            black_tx_m_read.address
			black_tx_m_read_waitrequest                      => black_tx_m_read_waitrequest,                                  --                                           .waitrequest
			black_tx_m_read_read                             => black_tx_m_read_read,                                         --                                           .read
			black_tx_m_read_readdata                         => black_tx_m_read_readdata,                                     --                                           .readdata
			black_tx_m_read_readdatavalid                    => black_tx_m_read_readdatavalid,                                --                                           .readdatavalid
			nios2_qsys_0_data_master_address                 => nios2_qsys_0_data_master_address,                             --                   nios2_qsys_0_data_master.address
			nios2_qsys_0_data_master_waitrequest             => nios2_qsys_0_data_master_waitrequest,                         --                                           .waitrequest
			nios2_qsys_0_data_master_byteenable              => nios2_qsys_0_data_master_byteenable,                          --                                           .byteenable
			nios2_qsys_0_data_master_read                    => nios2_qsys_0_data_master_read,                                --                                           .read
			nios2_qsys_0_data_master_readdata                => nios2_qsys_0_data_master_readdata,                            --                                           .readdata
			nios2_qsys_0_data_master_write                   => nios2_qsys_0_data_master_write,                               --                                           .write
			nios2_qsys_0_data_master_writedata               => nios2_qsys_0_data_master_writedata,                           --                                           .writedata
			nios2_qsys_0_data_master_debugaccess             => nios2_qsys_0_data_master_debugaccess,                         --                                           .debugaccess
			nios2_qsys_0_instruction_master_address          => nios2_qsys_0_instruction_master_address,                      --            nios2_qsys_0_instruction_master.address
			nios2_qsys_0_instruction_master_waitrequest      => nios2_qsys_0_instruction_master_waitrequest,                  --                                           .waitrequest
			nios2_qsys_0_instruction_master_read             => nios2_qsys_0_instruction_master_read,                         --                                           .read
			nios2_qsys_0_instruction_master_readdata         => nios2_qsys_0_instruction_master_readdata,                     --                                           .readdata
			red_rx_descriptor_read_address                   => red_rx_descriptor_read_address,                               --                     red_rx_descriptor_read.address
			red_rx_descriptor_read_waitrequest               => red_rx_descriptor_read_waitrequest,                           --                                           .waitrequest
			red_rx_descriptor_read_read                      => red_rx_descriptor_read_read,                                  --                                           .read
			red_rx_descriptor_read_readdata                  => red_rx_descriptor_read_readdata,                              --                                           .readdata
			red_rx_descriptor_read_readdatavalid             => red_rx_descriptor_read_readdatavalid,                         --                                           .readdatavalid
			red_rx_descriptor_write_address                  => red_rx_descriptor_write_address,                              --                    red_rx_descriptor_write.address
			red_rx_descriptor_write_waitrequest              => red_rx_descriptor_write_waitrequest,                          --                                           .waitrequest
			red_rx_descriptor_write_write                    => red_rx_descriptor_write_write,                                --                                           .write
			red_rx_descriptor_write_writedata                => red_rx_descriptor_write_writedata,                            --                                           .writedata
			red_rx_m_write_address                           => red_rx_m_write_address,                                       --                             red_rx_m_write.address
			red_rx_m_write_waitrequest                       => red_rx_m_write_waitrequest,                                   --                                           .waitrequest
			red_rx_m_write_byteenable                        => red_rx_m_write_byteenable,                                    --                                           .byteenable
			red_rx_m_write_write                             => red_rx_m_write_write,                                         --                                           .write
			red_rx_m_write_writedata                         => red_rx_m_write_writedata,                                     --                                           .writedata
			red_tx_descriptor_read_address                   => red_tx_descriptor_read_address,                               --                     red_tx_descriptor_read.address
			red_tx_descriptor_read_waitrequest               => red_tx_descriptor_read_waitrequest,                           --                                           .waitrequest
			red_tx_descriptor_read_read                      => red_tx_descriptor_read_read,                                  --                                           .read
			red_tx_descriptor_read_readdata                  => red_tx_descriptor_read_readdata,                              --                                           .readdata
			red_tx_descriptor_read_readdatavalid             => red_tx_descriptor_read_readdatavalid,                         --                                           .readdatavalid
			red_tx_descriptor_write_address                  => red_tx_descriptor_write_address,                              --                    red_tx_descriptor_write.address
			red_tx_descriptor_write_waitrequest              => red_tx_descriptor_write_waitrequest,                          --                                           .waitrequest
			red_tx_descriptor_write_write                    => red_tx_descriptor_write_write,                                --                                           .write
			red_tx_descriptor_write_writedata                => red_tx_descriptor_write_writedata,                            --                                           .writedata
			red_tx_m_read_address                            => red_tx_m_read_address,                                        --                              red_tx_m_read.address
			red_tx_m_read_waitrequest                        => red_tx_m_read_waitrequest,                                    --                                           .waitrequest
			red_tx_m_read_read                               => red_tx_m_read_read,                                           --                                           .read
			red_tx_m_read_readdata                           => red_tx_m_read_readdata,                                       --                                           .readdata
			red_tx_m_read_readdatavalid                      => red_tx_m_read_readdatavalid,                                  --                                           .readdatavalid
			ted_decryptor_read_master_address                => ted_decryptor_read_master_address,                            --                  ted_decryptor_read_master.address
			ted_decryptor_read_master_waitrequest            => ted_decryptor_read_master_waitrequest,                        --                                           .waitrequest
			ted_decryptor_read_master_read                   => ted_decryptor_read_master_read,                               --                                           .read
			ted_decryptor_read_master_readdata               => ted_decryptor_read_master_readdata,                           --                                           .readdata
			ted_decryptor_write_master_address               => ted_decryptor_write_master_address,                           --                 ted_decryptor_write_master.address
			ted_decryptor_write_master_waitrequest           => ted_decryptor_write_master_waitrequest,                       --                                           .waitrequest
			ted_decryptor_write_master_write                 => ted_decryptor_write_master_write,                             --                                           .write
			ted_decryptor_write_master_writedata             => ted_decryptor_write_master_writedata,                         --                                           .writedata
			ted_encryptor_read_master_address                => ted_encryptor_read_master_address,                            --                  ted_encryptor_read_master.address
			ted_encryptor_read_master_waitrequest            => ted_encryptor_read_master_waitrequest,                        --                                           .waitrequest
			ted_encryptor_read_master_read                   => ted_encryptor_read_master_read,                               --                                           .read
			ted_encryptor_read_master_readdata               => ted_encryptor_read_master_readdata,                           --                                           .readdata
			ted_encryptor_write_master_address               => ted_encryptor_write_master_address,                           --                 ted_encryptor_write_master.address
			ted_encryptor_write_master_waitrequest           => ted_encryptor_write_master_waitrequest,                       --                                           .waitrequest
			ted_encryptor_write_master_write                 => ted_encryptor_write_master_write,                             --                                           .write
			ted_encryptor_write_master_writedata             => ted_encryptor_write_master_writedata,                         --                                           .writedata
			black_interface_control_port_address             => mm_interconnect_0_black_interface_control_port_address,       --               black_interface_control_port.address
			black_interface_control_port_write               => mm_interconnect_0_black_interface_control_port_write,         --                                           .write
			black_interface_control_port_read                => mm_interconnect_0_black_interface_control_port_read,          --                                           .read
			black_interface_control_port_readdata            => mm_interconnect_0_black_interface_control_port_readdata,      --                                           .readdata
			black_interface_control_port_writedata           => mm_interconnect_0_black_interface_control_port_writedata,     --                                           .writedata
			black_interface_control_port_waitrequest         => mm_interconnect_0_black_interface_control_port_waitrequest,   --                                           .waitrequest
			black_rx_csr_address                             => mm_interconnect_0_black_rx_csr_address,                       --                               black_rx_csr.address
			black_rx_csr_write                               => mm_interconnect_0_black_rx_csr_write,                         --                                           .write
			black_rx_csr_read                                => mm_interconnect_0_black_rx_csr_read,                          --                                           .read
			black_rx_csr_readdata                            => mm_interconnect_0_black_rx_csr_readdata,                      --                                           .readdata
			black_rx_csr_writedata                           => mm_interconnect_0_black_rx_csr_writedata,                     --                                           .writedata
			black_rx_csr_chipselect                          => mm_interconnect_0_black_rx_csr_chipselect,                    --                                           .chipselect
			black_to_red_memory_s1_address                   => mm_interconnect_0_black_to_red_memory_s1_address,             --                     black_to_red_memory_s1.address
			black_to_red_memory_s1_write                     => mm_interconnect_0_black_to_red_memory_s1_write,               --                                           .write
			black_to_red_memory_s1_readdata                  => mm_interconnect_0_black_to_red_memory_s1_readdata,            --                                           .readdata
			black_to_red_memory_s1_writedata                 => mm_interconnect_0_black_to_red_memory_s1_writedata,           --                                           .writedata
			black_to_red_memory_s1_byteenable                => mm_interconnect_0_black_to_red_memory_s1_byteenable,          --                                           .byteenable
			black_to_red_memory_s1_chipselect                => mm_interconnect_0_black_to_red_memory_s1_chipselect,          --                                           .chipselect
			black_to_red_memory_s1_clken                     => mm_interconnect_0_black_to_red_memory_s1_clken,               --                                           .clken
			black_tx_csr_address                             => mm_interconnect_0_black_tx_csr_address,                       --                               black_tx_csr.address
			black_tx_csr_write                               => mm_interconnect_0_black_tx_csr_write,                         --                                           .write
			black_tx_csr_read                                => mm_interconnect_0_black_tx_csr_read,                          --                                           .read
			black_tx_csr_readdata                            => mm_interconnect_0_black_tx_csr_readdata,                      --                                           .readdata
			black_tx_csr_writedata                           => mm_interconnect_0_black_tx_csr_writedata,                     --                                           .writedata
			black_tx_csr_chipselect                          => mm_interconnect_0_black_tx_csr_chipselect,                    --                                           .chipselect
			descriptor_mem_s1_address                        => mm_interconnect_0_descriptor_mem_s1_address,                  --                          descriptor_mem_s1.address
			descriptor_mem_s1_write                          => mm_interconnect_0_descriptor_mem_s1_write,                    --                                           .write
			descriptor_mem_s1_readdata                       => mm_interconnect_0_descriptor_mem_s1_readdata,                 --                                           .readdata
			descriptor_mem_s1_writedata                      => mm_interconnect_0_descriptor_mem_s1_writedata,                --                                           .writedata
			descriptor_mem_s1_byteenable                     => mm_interconnect_0_descriptor_mem_s1_byteenable,               --                                           .byteenable
			descriptor_mem_s1_chipselect                     => mm_interconnect_0_descriptor_mem_s1_chipselect,               --                                           .chipselect
			descriptor_mem_s1_clken                          => mm_interconnect_0_descriptor_mem_s1_clken,                    --                                           .clken
			heap_stack_s1_address                            => mm_interconnect_0_heap_stack_s1_address,                      --                              heap_stack_s1.address
			heap_stack_s1_write                              => mm_interconnect_0_heap_stack_s1_write,                        --                                           .write
			heap_stack_s1_readdata                           => mm_interconnect_0_heap_stack_s1_readdata,                     --                                           .readdata
			heap_stack_s1_writedata                          => mm_interconnect_0_heap_stack_s1_writedata,                    --                                           .writedata
			heap_stack_s1_byteenable                         => mm_interconnect_0_heap_stack_s1_byteenable,                   --                                           .byteenable
			heap_stack_s1_chipselect                         => mm_interconnect_0_heap_stack_s1_chipselect,                   --                                           .chipselect
			heap_stack_s1_clken                              => mm_interconnect_0_heap_stack_s1_clken,                        --                                           .clken
			hex_avalon_slave_0_write                         => mm_interconnect_0_hex_avalon_slave_0_write,                   --                         hex_avalon_slave_0.write
			hex_avalon_slave_0_read                          => mm_interconnect_0_hex_avalon_slave_0_read,                    --                                           .read
			hex_avalon_slave_0_readdata                      => mm_interconnect_0_hex_avalon_slave_0_readdata,                --                                           .readdata
			hex_avalon_slave_0_writedata                     => mm_interconnect_0_hex_avalon_slave_0_writedata,               --                                           .writedata
			hex_avalon_slave_0_byteenable                    => mm_interconnect_0_hex_avalon_slave_0_byteenable,              --                                           .byteenable
			hex_avalon_slave_0_chipselect                    => mm_interconnect_0_hex_avalon_slave_0_chipselect,              --                                           .chipselect
			input_port_s1_address                            => mm_interconnect_0_input_port_s1_address,                      --                              input_port_s1.address
			input_port_s1_readdata                           => mm_interconnect_0_input_port_s1_readdata,                     --                                           .readdata
			instruction_memory_s1_address                    => mm_interconnect_0_instruction_memory_s1_address,              --                      instruction_memory_s1.address
			instruction_memory_s1_write                      => mm_interconnect_0_instruction_memory_s1_write,                --                                           .write
			instruction_memory_s1_readdata                   => mm_interconnect_0_instruction_memory_s1_readdata,             --                                           .readdata
			instruction_memory_s1_writedata                  => mm_interconnect_0_instruction_memory_s1_writedata,            --                                           .writedata
			instruction_memory_s1_byteenable                 => mm_interconnect_0_instruction_memory_s1_byteenable,           --                                           .byteenable
			instruction_memory_s1_chipselect                 => mm_interconnect_0_instruction_memory_s1_chipselect,           --                                           .chipselect
			instruction_memory_s1_clken                      => mm_interconnect_0_instruction_memory_s1_clken,                --                                           .clken
			jtag_uart_avalon_jtag_slave_address              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,        --                jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,          --                                           .write
			jtag_uart_avalon_jtag_slave_read                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,           --                                           .read
			jtag_uart_avalon_jtag_slave_readdata             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,       --                                           .readdata
			jtag_uart_avalon_jtag_slave_writedata            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,      --                                           .writedata
			jtag_uart_avalon_jtag_slave_waitrequest          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,    --                                           .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,     --                                           .chipselect
			lcd_avalon_lcd_slave_address                     => mm_interconnect_0_lcd_avalon_lcd_slave_address,               --                       lcd_avalon_lcd_slave.address
			lcd_avalon_lcd_slave_write                       => mm_interconnect_0_lcd_avalon_lcd_slave_write,                 --                                           .write
			lcd_avalon_lcd_slave_read                        => mm_interconnect_0_lcd_avalon_lcd_slave_read,                  --                                           .read
			lcd_avalon_lcd_slave_readdata                    => mm_interconnect_0_lcd_avalon_lcd_slave_readdata,              --                                           .readdata
			lcd_avalon_lcd_slave_writedata                   => mm_interconnect_0_lcd_avalon_lcd_slave_writedata,             --                                           .writedata
			lcd_avalon_lcd_slave_waitrequest                 => mm_interconnect_0_lcd_avalon_lcd_slave_waitrequest,           --                                           .waitrequest
			lcd_avalon_lcd_slave_chipselect                  => mm_interconnect_0_lcd_avalon_lcd_slave_chipselect,            --                                           .chipselect
			lcd_clk_pll_slave_address                        => mm_interconnect_0_lcd_clk_pll_slave_address,                  --                          lcd_clk_pll_slave.address
			lcd_clk_pll_slave_write                          => mm_interconnect_0_lcd_clk_pll_slave_write,                    --                                           .write
			lcd_clk_pll_slave_read                           => mm_interconnect_0_lcd_clk_pll_slave_read,                     --                                           .read
			lcd_clk_pll_slave_readdata                       => mm_interconnect_0_lcd_clk_pll_slave_readdata,                 --                                           .readdata
			lcd_clk_pll_slave_writedata                      => mm_interconnect_0_lcd_clk_pll_slave_writedata,                --                                           .writedata
			nios2_qsys_0_jtag_debug_module_address           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --             nios2_qsys_0_jtag_debug_module.address
			nios2_qsys_0_jtag_debug_module_write             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                                           .write
			nios2_qsys_0_jtag_debug_module_read              => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                                           .read
			nios2_qsys_0_jtag_debug_module_readdata          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                                           .readdata
			nios2_qsys_0_jtag_debug_module_writedata         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                                           .writedata
			nios2_qsys_0_jtag_debug_module_byteenable        => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                                           .byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                                           .waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess       => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                                           .debugaccess
			output_port_s1_address                           => mm_interconnect_0_output_port_s1_address,                     --                             output_port_s1.address
			output_port_s1_write                             => mm_interconnect_0_output_port_s1_write,                       --                                           .write
			output_port_s1_readdata                          => mm_interconnect_0_output_port_s1_readdata,                    --                                           .readdata
			output_port_s1_writedata                         => mm_interconnect_0_output_port_s1_writedata,                   --                                           .writedata
			output_port_s1_chipselect                        => mm_interconnect_0_output_port_s1_chipselect,                  --                                           .chipselect
			red_interface_control_port_address               => mm_interconnect_0_red_interface_control_port_address,         --                 red_interface_control_port.address
			red_interface_control_port_write                 => mm_interconnect_0_red_interface_control_port_write,           --                                           .write
			red_interface_control_port_read                  => mm_interconnect_0_red_interface_control_port_read,            --                                           .read
			red_interface_control_port_readdata              => mm_interconnect_0_red_interface_control_port_readdata,        --                                           .readdata
			red_interface_control_port_writedata             => mm_interconnect_0_red_interface_control_port_writedata,       --                                           .writedata
			red_interface_control_port_waitrequest           => mm_interconnect_0_red_interface_control_port_waitrequest,     --                                           .waitrequest
			red_rx_csr_address                               => mm_interconnect_0_red_rx_csr_address,                         --                                 red_rx_csr.address
			red_rx_csr_write                                 => mm_interconnect_0_red_rx_csr_write,                           --                                           .write
			red_rx_csr_read                                  => mm_interconnect_0_red_rx_csr_read,                            --                                           .read
			red_rx_csr_readdata                              => mm_interconnect_0_red_rx_csr_readdata,                        --                                           .readdata
			red_rx_csr_writedata                             => mm_interconnect_0_red_rx_csr_writedata,                       --                                           .writedata
			red_rx_csr_chipselect                            => mm_interconnect_0_red_rx_csr_chipselect,                      --                                           .chipselect
			red_to_black_memory_s1_address                   => mm_interconnect_0_red_to_black_memory_s1_address,             --                     red_to_black_memory_s1.address
			red_to_black_memory_s1_write                     => mm_interconnect_0_red_to_black_memory_s1_write,               --                                           .write
			red_to_black_memory_s1_readdata                  => mm_interconnect_0_red_to_black_memory_s1_readdata,            --                                           .readdata
			red_to_black_memory_s1_writedata                 => mm_interconnect_0_red_to_black_memory_s1_writedata,           --                                           .writedata
			red_to_black_memory_s1_byteenable                => mm_interconnect_0_red_to_black_memory_s1_byteenable,          --                                           .byteenable
			red_to_black_memory_s1_chipselect                => mm_interconnect_0_red_to_black_memory_s1_chipselect,          --                                           .chipselect
			red_to_black_memory_s1_clken                     => mm_interconnect_0_red_to_black_memory_s1_clken,               --                                           .clken
			red_tx_csr_address                               => mm_interconnect_0_red_tx_csr_address,                         --                                 red_tx_csr.address
			red_tx_csr_write                                 => mm_interconnect_0_red_tx_csr_write,                           --                                           .write
			red_tx_csr_read                                  => mm_interconnect_0_red_tx_csr_read,                            --                                           .read
			red_tx_csr_readdata                              => mm_interconnect_0_red_tx_csr_readdata,                        --                                           .readdata
			red_tx_csr_writedata                             => mm_interconnect_0_red_tx_csr_writedata,                       --                                           .writedata
			red_tx_csr_chipselect                            => mm_interconnect_0_red_tx_csr_chipselect,                      --                                           .chipselect
			system_id_control_slave_address                  => mm_interconnect_0_system_id_control_slave_address,            --                    system_id_control_slave.address
			system_id_control_slave_readdata                 => mm_interconnect_0_system_id_control_slave_readdata,           --                                           .readdata
			system_timer_s1_address                          => mm_interconnect_0_system_timer_s1_address,                    --                            system_timer_s1.address
			system_timer_s1_write                            => mm_interconnect_0_system_timer_s1_write,                      --                                           .write
			system_timer_s1_readdata                         => mm_interconnect_0_system_timer_s1_readdata,                   --                                           .readdata
			system_timer_s1_writedata                        => mm_interconnect_0_system_timer_s1_writedata,                  --                                           .writedata
			system_timer_s1_chipselect                       => mm_interconnect_0_system_timer_s1_chipselect,                 --                                           .chipselect
			ted_decryptor_csr_address                        => mm_interconnect_0_ted_decryptor_csr_address,                  --                          ted_decryptor_csr.address
			ted_decryptor_csr_write                          => mm_interconnect_0_ted_decryptor_csr_write,                    --                                           .write
			ted_decryptor_csr_readdata                       => mm_interconnect_0_ted_decryptor_csr_readdata,                 --                                           .readdata
			ted_decryptor_csr_writedata                      => mm_interconnect_0_ted_decryptor_csr_writedata,                --                                           .writedata
			ted_encryptor_csr_address                        => mm_interconnect_0_ted_encryptor_csr_address,                  --                          ted_encryptor_csr.address
			ted_encryptor_csr_write                          => mm_interconnect_0_ted_encryptor_csr_write,                    --                                           .write
			ted_encryptor_csr_readdata                       => mm_interconnect_0_ted_encryptor_csr_readdata,                 --                                           .readdata
			ted_encryptor_csr_writedata                      => mm_interconnect_0_ted_encryptor_csr_writedata                 --                                           .writedata
		);

	irq_mapper : component TEDv3_architecture_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,       -- receiver5.irq
			sender_irq    => nios2_qsys_0_d_irq_irq          --    sender.irq
		);

	avalon_st_adapter : component TEDv3_architecture_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 1,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                               -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,        -- in_rst_0.reset
			in_0_data           => black_tx_out_data,                     --     in_0.data
			in_0_valid          => black_tx_out_valid,                    --         .valid
			in_0_ready          => black_tx_out_ready,                    --         .ready
			in_0_startofpacket  => black_tx_out_startofpacket,            --         .startofpacket
			in_0_endofpacket    => black_tx_out_endofpacket,              --         .endofpacket
			in_0_empty          => black_tx_out_empty,                    --         .empty
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	avalon_st_adapter_001 : component TEDv3_architecture_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 1,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                                   -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,            -- in_rst_0.reset
			in_0_data           => red_tx_out_data,                           --     in_0.data
			in_0_valid          => red_tx_out_valid,                          --         .valid
			in_0_ready          => red_tx_out_ready,                          --         .ready
			in_0_startofpacket  => red_tx_out_startofpacket,                  --         .startofpacket
			in_0_endofpacket    => red_tx_out_endofpacket,                    --         .endofpacket
			in_0_empty          => red_tx_out_empty,                          --         .empty
			out_0_data          => avalon_st_adapter_001_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_001_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_001_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_001_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_001_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_001_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_001_out_0_error          --         .error
		);

	avalon_st_adapter_002 : component TEDv3_architecture_avalon_st_adapter_002
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                                   -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,            -- in_rst_0.reset
			in_0_data           => black_interface_receive_data,              --     in_0.data
			in_0_valid          => black_interface_receive_valid,             --         .valid
			in_0_ready          => black_interface_receive_ready,             --         .ready
			in_0_startofpacket  => black_interface_receive_startofpacket,     --         .startofpacket
			in_0_endofpacket    => black_interface_receive_endofpacket,       --         .endofpacket
			in_0_empty          => black_interface_receive_empty,             --         .empty
			in_0_error          => black_interface_receive_error,             --         .error
			out_0_data          => avalon_st_adapter_002_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_002_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_002_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_002_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_002_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_002_out_0_empty          --         .empty
		);

	avalon_st_adapter_003 : component TEDv3_architecture_avalon_st_adapter_002
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                                   -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,            -- in_rst_0.reset
			in_0_data           => red_interface_receive_data,                --     in_0.data
			in_0_valid          => red_interface_receive_valid,               --         .valid
			in_0_ready          => red_interface_receive_ready,               --         .ready
			in_0_startofpacket  => red_interface_receive_startofpacket,       --         .startofpacket
			in_0_endofpacket    => red_interface_receive_endofpacket,         --         .endofpacket
			in_0_empty          => red_interface_receive_empty,               --         .empty
			in_0_error          => red_interface_receive_error,               --         .error
			out_0_data          => avalon_st_adapter_003_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_003_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_003_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_003_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_003_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_003_out_0_empty          --         .empty
		);

	rst_controller : component tedv3_architecture_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clk_clk,                                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,         --          .reset_req
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_001 : component tedv3_architecture_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => lcd_clk_c0_clk,                             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_output_port_s1_write_ports_inv <= not mm_interconnect_0_output_port_s1_write;

	mm_interconnect_0_system_timer_s1_write_ports_inv <= not mm_interconnect_0_system_timer_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of TEDv3_architecture
