
module TEDv3_architecture (
	black_interface_mac_mdio_connection_mdc,
	black_interface_mac_mdio_connection_mdio_in,
	black_interface_mac_mdio_connection_mdio_out,
	black_interface_mac_mdio_connection_mdio_oen,
	black_interface_mac_misc_connection_xon_gen,
	black_interface_mac_misc_connection_xoff_gen,
	black_interface_mac_misc_connection_ff_tx_crc_fwd,
	black_interface_mac_misc_connection_ff_tx_septy,
	black_interface_mac_misc_connection_tx_ff_uflow,
	black_interface_mac_misc_connection_ff_tx_a_full,
	black_interface_mac_misc_connection_ff_tx_a_empty,
	black_interface_mac_misc_connection_rx_err_stat,
	black_interface_mac_misc_connection_rx_frm_type,
	black_interface_mac_misc_connection_ff_rx_dsav,
	black_interface_mac_misc_connection_ff_rx_a_full,
	black_interface_mac_misc_connection_ff_rx_a_empty,
	black_interface_mac_rgmii_connection_rgmii_in,
	black_interface_mac_rgmii_connection_rgmii_out,
	black_interface_mac_rgmii_connection_rx_control,
	black_interface_mac_rgmii_connection_tx_control,
	black_interface_mac_status_connection_set_10,
	black_interface_mac_status_connection_set_1000,
	black_interface_mac_status_connection_eth_mode,
	black_interface_mac_status_connection_ena_10,
	black_interface_pcs_mac_rx_clock_connection_clk,
	black_interface_pcs_mac_tx_clock_connection_clk,
	clk_clk,
	hex_conduit_hex_conduit,
	input_port_external_connection_export,
	lcd_clk_areset_conduit_export,
	lcd_clk_locked_conduit_export,
	lcd_clk_phasedone_conduit_export,
	lcd_external_interface_DATA,
	lcd_external_interface_ON,
	lcd_external_interface_BLON,
	lcd_external_interface_EN,
	lcd_external_interface_RS,
	lcd_external_interface_RW,
	output_port_external_connection_export,
	red_interface_mac_mdio_connection_mdc,
	red_interface_mac_mdio_connection_mdio_in,
	red_interface_mac_mdio_connection_mdio_out,
	red_interface_mac_mdio_connection_mdio_oen,
	red_interface_mac_misc_connection_xon_gen,
	red_interface_mac_misc_connection_xoff_gen,
	red_interface_mac_misc_connection_ff_tx_crc_fwd,
	red_interface_mac_misc_connection_ff_tx_septy,
	red_interface_mac_misc_connection_tx_ff_uflow,
	red_interface_mac_misc_connection_ff_tx_a_full,
	red_interface_mac_misc_connection_ff_tx_a_empty,
	red_interface_mac_misc_connection_rx_err_stat,
	red_interface_mac_misc_connection_rx_frm_type,
	red_interface_mac_misc_connection_ff_rx_dsav,
	red_interface_mac_misc_connection_ff_rx_a_full,
	red_interface_mac_misc_connection_ff_rx_a_empty,
	red_interface_mac_rgmii_connection_rgmii_in,
	red_interface_mac_rgmii_connection_rgmii_out,
	red_interface_mac_rgmii_connection_rx_control,
	red_interface_mac_rgmii_connection_tx_control,
	red_interface_mac_status_connection_set_10,
	red_interface_mac_status_connection_set_1000,
	red_interface_mac_status_connection_eth_mode,
	red_interface_mac_status_connection_ena_10,
	red_interface_pcs_mac_rx_clock_connection_clk,
	red_interface_pcs_mac_tx_clock_connection_clk,
	reset_reset_n);	

	output		black_interface_mac_mdio_connection_mdc;
	input		black_interface_mac_mdio_connection_mdio_in;
	output		black_interface_mac_mdio_connection_mdio_out;
	output		black_interface_mac_mdio_connection_mdio_oen;
	input		black_interface_mac_misc_connection_xon_gen;
	input		black_interface_mac_misc_connection_xoff_gen;
	input		black_interface_mac_misc_connection_ff_tx_crc_fwd;
	output		black_interface_mac_misc_connection_ff_tx_septy;
	output		black_interface_mac_misc_connection_tx_ff_uflow;
	output		black_interface_mac_misc_connection_ff_tx_a_full;
	output		black_interface_mac_misc_connection_ff_tx_a_empty;
	output	[17:0]	black_interface_mac_misc_connection_rx_err_stat;
	output	[3:0]	black_interface_mac_misc_connection_rx_frm_type;
	output		black_interface_mac_misc_connection_ff_rx_dsav;
	output		black_interface_mac_misc_connection_ff_rx_a_full;
	output		black_interface_mac_misc_connection_ff_rx_a_empty;
	input	[3:0]	black_interface_mac_rgmii_connection_rgmii_in;
	output	[3:0]	black_interface_mac_rgmii_connection_rgmii_out;
	input		black_interface_mac_rgmii_connection_rx_control;
	output		black_interface_mac_rgmii_connection_tx_control;
	input		black_interface_mac_status_connection_set_10;
	input		black_interface_mac_status_connection_set_1000;
	output		black_interface_mac_status_connection_eth_mode;
	output		black_interface_mac_status_connection_ena_10;
	input		black_interface_pcs_mac_rx_clock_connection_clk;
	input		black_interface_pcs_mac_tx_clock_connection_clk;
	input		clk_clk;
	output	[31:0]	hex_conduit_hex_conduit;
	input	[31:0]	input_port_external_connection_export;
	input		lcd_clk_areset_conduit_export;
	output		lcd_clk_locked_conduit_export;
	output		lcd_clk_phasedone_conduit_export;
	inout	[7:0]	lcd_external_interface_DATA;
	output		lcd_external_interface_ON;
	output		lcd_external_interface_BLON;
	output		lcd_external_interface_EN;
	output		lcd_external_interface_RS;
	output		lcd_external_interface_RW;
	output	[31:0]	output_port_external_connection_export;
	output		red_interface_mac_mdio_connection_mdc;
	input		red_interface_mac_mdio_connection_mdio_in;
	output		red_interface_mac_mdio_connection_mdio_out;
	output		red_interface_mac_mdio_connection_mdio_oen;
	input		red_interface_mac_misc_connection_xon_gen;
	input		red_interface_mac_misc_connection_xoff_gen;
	input		red_interface_mac_misc_connection_ff_tx_crc_fwd;
	output		red_interface_mac_misc_connection_ff_tx_septy;
	output		red_interface_mac_misc_connection_tx_ff_uflow;
	output		red_interface_mac_misc_connection_ff_tx_a_full;
	output		red_interface_mac_misc_connection_ff_tx_a_empty;
	output	[17:0]	red_interface_mac_misc_connection_rx_err_stat;
	output	[3:0]	red_interface_mac_misc_connection_rx_frm_type;
	output		red_interface_mac_misc_connection_ff_rx_dsav;
	output		red_interface_mac_misc_connection_ff_rx_a_full;
	output		red_interface_mac_misc_connection_ff_rx_a_empty;
	input	[3:0]	red_interface_mac_rgmii_connection_rgmii_in;
	output	[3:0]	red_interface_mac_rgmii_connection_rgmii_out;
	input		red_interface_mac_rgmii_connection_rx_control;
	output		red_interface_mac_rgmii_connection_tx_control;
	input		red_interface_mac_status_connection_set_10;
	input		red_interface_mac_status_connection_set_1000;
	output		red_interface_mac_status_connection_eth_mode;
	output		red_interface_mac_status_connection_ena_10;
	input		red_interface_pcs_mac_rx_clock_connection_clk;
	input		red_interface_pcs_mac_tx_clock_connection_clk;
	input		reset_reset_n;
endmodule
