// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1.1
// ALTERA_TIMESTAMP:Tue Jan 20 08:33:55 PST 2015
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k1CowpfWzXzbz3BsY6XNPBIjVlw9XyrNhhstU2pPR4yGJUHsP4JwRcUde3QRIV/1
x78NzrHC1ESvIAPvxSGfnpcM1OuJsHi9ro6Z+aQceJQYwWpm3bXCER1/muSjTdUf
5V19Qf1ycMJevn1k0hLFytBG4Gvhue5eXZxDePNUA9c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29408)
Pb3eTmD5HJsiV9xbJKJ3kycEZrma7bzjmyjyOqAFI276AlWw8/CMal7OuFmR5q7o
sWV/TBgH+ApZFUsuBH1Nkyf3dEu9TYYedlmfE0o33i/6+nf+IedUt0Dmcc7b2Bxz
G62CsL0wNG3AsMG6Khax0Km+Z+KBAyUNmDl9RURJxRfPOZav7CYIqtTygkubvoWV
wwzNAtWhQYZk/Ey9HicLa+MhTcUb2VUOwrIz/XDNgXuk0VbzXYZ83JipVJPQIasR
e8z6EGIwaIhFjYwJCyl3VyS2p3HSMKI0DJZUWowQUjiHzUTvmPO15jNtuwYgCs0r
Slgz99Gl3KQa7ujvRLddlwBTFXaQF7p3bk4Vdm5XsUBMsaWM/Gd603yQ7h9UPNWD
gOVdEbZSHPzDsZZRMrfY6a6x11PMMGfLaNXZbLlEFJtw8RUXDJ0ix/2sLkpw59xR
hLGz9eb8SaZhwkcAl/6HQVPMYsVjon0zv624ZAfrdbU369WGdy/Gxnu0wrno8GKU
CVgnyHGZ3Sq7LOGEJ1ZhZ2HaM0iCuCslDtlYwqpF1Q1KyotusXCFzJ1gpXRvz+hc
lwY8ZS4eb7fEAClkRhvM01TV3FKmIEWls3yBFeglUQqsyB2OHvoc5UqB34FuV+Ie
XuXiZp+WpLifTM6cX+wmWKD4E7oSdqvvBT/2FnF8ZUnmnlsP0MxnLbKTAKc8YOdt
I3mWeJ5QldomslcdVpeCixU2TgV/lkG27yEqHiCTBo10ukzth6cGzPEJHeanYALF
l51Zxw+JTp9ieqtugh93JvKW854C1yLB8UzqUGy/5o9w91W8nl8jc6244KhUzQG0
PTmdtZrI6dvjOLF0SahemFFHBqeceSk7wh4O0Rae3qAm5UkUhGdaVzlIrLFJspTc
hgI/gHxJRuxSydN8uWMjkvy+t8P9kZoJ/1dA22ouzSuX/rLlSqdRiOwtT+sFrnzH
31xdKakYtxciP8MbATm8zNzz9NnVXvbC1Gksb0aNismBhU5gv8vkWqP+epylZPl6
l19hJ3Od+z5iGuDw5uXhd3HSsLYZIyM+ck/KuuSjRC/FjbJd6Y7d3A9j8SmBfjcU
KAJ5Tzd7EUhEz2AVD1nyHkROuO1k0ExGA7igP6uZmE1WKwMV9EepCF+bUT5F+tfo
BAk4m3BrA4OLVsAazNWGDrKmDnmkLPsDq1r3nitu77FrYFmlX2/iCgennS8Y9E8l
efd5gg5iKIRSpLE+29eOusH5fGcF8VgTKrk76aJTwQ3Ny7CFT3GcsvG5b+KMjWGX
4jUYHTKsFYHKZ+NCQdmDULpjgXCgKKBdF8pdp2TAa5gljUSSt4i9qMR3zpv4bFVj
VDb61VYceJ6EV/q4wb/cUrkG6orqixFth6DbhsQG3dN8Lc4sGOHMzJOn+j7CORgY
/bXkT9NHuDksyhW13F5mImSHVeG9g1iBSLLq3sBKj4wfkT6nqmbbyeRgowsozysS
QDTTaDbmW9OEmjQtAo0qAY8QKN6Hy9JijmM73wPTcqi8M+zZRUP1S77ClyGR9Hk+
Od5BTOeKXolO1wGYuOUTbbRF6Ohz1H8m43Y0IEfU4glujsMo5xJTg21+NwNAD7jZ
jeHCHTmOnQiQaRb9srodnbGf0N3xvQ7ikR1JeAZYA9XorGoc+/HXMbPe0Y+WUBiH
1GHGwu5zm1auiNXMDlYF5oMsKgaJ/N/N+CdF3vZZWfsAdtKd919DZiVytArOoPir
G3xJ96jYkzp9tS5H9x5d4pJN0YcHT0zDHMflUNgSE7whmVB2R6k5zmRYhCmhB0CS
ASeirZDPAOMQtUUnay5TAiAG773+O202DcyLTXtkkb1mIH15R9ux6ZsNPZUgAAnL
1eDdJF2sGCaOMRFhX7XGM/T1m7DhEs9oZGBfqyiVo5dF/hYxDzXwlaI3yds7qTN9
3CEWRxNBTKcWRwGXkN7JVbf1TAdYHrq7jKFzv6mXCLpi+4cZN0m7B9xsXx6IhxsP
v7cHq3S3d2n4VfCCfuVWLXEcef7ll+nPa6Mic3S+yDJU4Mt/TGM10U+zYwfx2zb0
z0JFlC8SaOKGiHRb9/z+yn6tBulh5KWdXCQcK5ERZb+E/pjzxfzZl/i2HkE+U0F4
ShED+9dW8kJzVSRwT2L8FHBkariMkZJUJa39cRiBGyYewo9ZU/Pe1SOTK/A1HtVp
I7cWzzEGWHJnAIKoxDTVE0KuO1gcLfI9NxJUMwmsSZb1frDkv7B+rOMpHWTVoAiB
dGn6w/XFVt6fcscMMrUo8pGqWlukzpzzzuvhUQtRWK32WhwiZGKyY76Wb3XEvD23
7Gff50tggXSqsd70GPIDYlMarmYNHWo9FJPf0r2IZ+Pu2nRSqN+pCv6uDhOaVq7L
cVl6LHcJ4vLdk4Lvwz89rSUnghBjeFdyKn2LxfBQZHgYlkgTb6dkCs75wxFfBNWy
/sVE49nflIOAguVyF8MaO5anjjKCtTm3VAXXGPeVXLzZcAO/87laLh/YxaBgU7W1
WpdUA5lyWCshp944buk4v7MqJQgBgmVE7hY0MGQ7QvVLcUsyzH2BLnwT+IPZn09M
0LqiW7r/jlNngpiI5/RlIcjwqntdBm492yi9AHrGUIpOWBPdEwHa4xXTUUA22W9P
Ec9lvDuWsId8m89EDC0BYOwP7RH/FaV+8EHgGxaLjfzOLawD40OTUiSjPodEtBtm
d2JgOY7kr05AKBx5MmndQKqxX+3oRR1MDTQkXMCShH7ltObXI0eJGzHR67LQeiE8
2Wx3QhLlLH2i7lpz1tnjnoL+k9Vx5Y+cwW5zznz9gmJfcKfr0emFjVRSM9ncpgeU
WzBIn8fzqLWfye6SiG+OsN7eBOybUMhGY6fZjG0p74wCW/GEMqS+Mh1ntS+QQ3bR
c8ijr27YrF2M7+UH7zOoeDtXUYaseOKjDIJIkW4zFe8J7813J9oSVsfNx1qYmF/E
RDRvDk+BdvoEhPH+tENhsYo7asUh28WN9EuSJ5uYEBCuHNGcZOVaBmTEtcs2L4+t
yV8MOn8gzBgnbyHFTXfStUZe0bl6+vwiy+f5j2KsYIckNrGqs4YGnQIEAR51e4he
28drxkw+Q7jGLCkWYnTXvSChDrsM5FZaG5fWVlQrVJKDWzLRUS3wscPu65RqtZoB
kXSyj3+V0EggT30R5RjDlflWQeo7ujTMDvNgqH0SZqYHj04fj6YbbS/Q0ZRoCYQt
N2SEPcdF0Pwj2ggMsV9+eDRETsmYqUtVlqkL20gOCEdn34H1JT0LqQdrStzBDDnt
SseSRECeW0gFUQIIGlLibYCJmxBE3XkxctrOM7qUNnzC3uRqhUKSHaTnnY3KFIaA
MU2rUFK5uuziaT5+Loc3TVEqKAY229/reO5+b1zj4iGrBZNLwUsF5muS4Z2A7e7F
Sb03JWTSBZ8hobcRCYYcUnh51X5VZ1NmWkfHWpzb9ZVNUhIIPd5LAVA1ezKjLphW
kossbOchOJvsm0cPwmGJHXPbgb8di9JjZuguNGiRpmG6mL9zFSCKeTJVs1ei34g5
HVasWRYYNLfw/WvvK7cP0uWGmTe8yENsq5KZiHug1T/h+2cEkpJ1CsnLb7cQnyTm
IUvkoCX8pf7WorwTfSgjB4TAlGPSVeEIOyNXeBqiPfub1IT7fCX7krwX5IOiWGzM
+ry2h/Gi+Ud9iFSqCorer3SC7dYjM6eyIdL/d2kd6uZgMS8Ce+KrIjXSUw98VpBd
3YbiYSygyAPn1VzKE0pBt+FoKYrFpRGKEEkW1RmLYVOiZYhEK7Fdzb3YpB8ZErhu
UFgiZzoTM3gOujykRncNtxaOhX9/+SP87vWVnG6y5k6Nm8DpScWHYpagQS8+Z3G1
IWV7n58N/GNtwJi5MxXh16FDvoIt4VRneW5TngiThH22XeCWrYPMY62Beh54/jyB
M7t3ii3n07DWlr9+3McDBIV7xbx5z+tbb+1NZv2BRXxAmjrAXq5d1jw6vBD7+UNp
ZIiw6qt/Tf0d4i+IVhV6PjN/ktjC5/Ny73IfkFDWtJNNOd/gtDBaRpVy9m4ppOVg
+eA3YwgarD1TynJA13M96fOHi/DKW9iSfe4f3pusD/IrXv9UeZBDa6+oTssS8RVY
rWZ2H9sWH+RxwTWaVMNDZqYRh4qfgIbygcFRwfF6hucM9Bp7KaMj8lgd0bn5g5I1
MVKYhDkPsQbacERZx/Qslk9RC9V7LLM24ad1UHoaH9UJnlXbm7gLBxYRhL3vfVDL
FWXI7j6gezdaqFgKAtbpxfuBSnWuLBmYwdo/U6GpjxcRO1pqf2uBimUryuNzAupF
pCoeyxT+8+HTTkka3gIsA7Aq4SWiICd7dYBD6hqpwg1MTzET5pt1vLFvfulf0744
5q211dgA9tHjavH6gLXrPzhFvHYtnMVuCMs/GCzeb2exVnayBsYJOor7PwBuRA3M
O16voY+if+zZvo+2R9ww1zB0F0mF2MzSMXjv5DZdM+C+gG/HRhuOHDFjGv72v19F
TsbYPZj+uRt5imXbtsb+lRfgUWl+Xsx4EdvZ0do9/JISEGdqvVtFNR4FNmyTj4ip
EoCz0behCkvP54Q2h8Au0o/jgTYnETM3lM6xse4sC2p6giUJS6gbGXsSM0wg0W/J
XdZcU444hMwtGlZiEduIsupkf0cANdOVKgODwGHhm63+/Ax5YgMRAZK+VA6jsPlT
o7o1tLg0H0ZkZiHwCe1jR2ELBxfS7WScLf8CgOGvBH3VQZHQWPzTzwIayx8UfJI/
qIFnYkvyxsUwBWgniz9cvPBO84ax/L6KbBVgklGV10mOsyYsCuzffMXhlXBsge9L
QGamjDGidnSUOgADFBd0SNx+syyrZ/BWV7D8oekiGrJ0cCIhma1XfurAisU1g/sE
i2sBbLL/NrOD/7kXdT6s4cJYcxP+U6EVTW3wWnt6xYt8JN/ZKSJYwoucaUU1HWdZ
Sc2sHoJcGYKj94Emr8qlr1nYxsM9vQcP+PNPBToe1iOaMsOD8/fBOEwC2MRO8RjE
bRgN6M+IvqUWWb4sviCPXWbrvvn03nWoM0QOOSJQcH7+Sib0tqewOmydMJp0vJhJ
pIDvdoN2gOaHYR7FTaIm9UKkBZupuGKseRzX0CJi6twZ7qfVvrzQrJsmyC3dWV0I
JEb0+651T8C/9NxapOhHGuG6cIM4B6DSd1UCUbZsWPnxaYfNsDX3NhQ8QEwK5x3t
9QXk5/vpIPvZcDgroDt4ki+jPHHusIHHLP9ymfetpGfNuUEf3hAstQ/7N7XKm2MK
dxp7G5ZNvdRF5q+1Gvi+S0KVUdaPf8BKwdUVf/5EfRdOxIbP4LaKlntpgQJf3bZi
HM2HGpSy9bhip2D7YhBL8JGZw5neE0JtcZm6NhjmOsgbSU5cmrO5iyV1LyGLY+Fo
Jjwy6UkAYL15GtJaB43LJpJlJnqtISKizWvzoSFud64PQz5nNopmccJ7Qq6MZ8ks
UXC7LbLyboq3viDHxpZd5fSlaCE7j7X6TrDVsQ+NHp9dFT3zcba/A6vqYNFYT6oe
ecq+ZrkcD3M/HXXIBZPv7qvi9FgLYSUV8tSHqHC9xZK8QTw99C/dByNxsW8dyuUe
dU0QMpm9m2NU6H7730YfC4D/c7CjbRgfwqjA5MDvOw3npJsxSlbmXDUso3GYyIJ3
dcQKSeZbxJek7aiA2/v+Yqr5lsrBqnSm5J/Ui5vNXUpAkbwGquG9qEH3SQlZwLxZ
1ftN3YZmCWWyJhUkeqkTXYecsSd01uLh4V6TgCHq1Ch+j/b8YonVdU5sRu+tuRcI
+Sp947LcTw5YEFBlPTFb6ycdb8Xm5mvVOZ3pYNdIuKQft8apI/6TGxXG4dS9BToA
FXGugwSjDm6lBMwe0uyrodLkGXx7oPT3+44Kc7qw8DCQsS6rfEoa+CnO6Z3Cogdc
ETuBq5Nu2uyseYTh7J1kxcmeMqcR5rCRgJKBB2aui6KmwaYSdOx1Sv/yUGvRLKPb
D50oHDHn0D3zFSipNmzY1QCceQphF4uGGN08N3GdnJIHibRYl6exOOif6CHiZn/I
cerZljKDEgauH+qJLkoqWOMepFP4ZZ1JHtdwan9tzvsVZF7VugAexiS+ax7MG4W9
m3Ms4VjErE9WRNZ2LLZkYln2yHAvsB4ULA1zsP2qyFDsPjXx/462EWeCfUd0RRQ2
cgTiTXkXUfaBxgMYHJCHS1lNDeAho8RxWei6+1Q4444RW1n+kcvxe68l5WPJDKjf
FqJsBznzjQvCvb63KJIcmbWVJ3NyGPIaifHqYsUx1644oSLijbzMbSiRUwp73mCL
aF9RMgTyrLRoUTKs1mh0gGwrxyGcQc5bWctvSznH2P5GkiXuV5JVOx1zpcMuVHwX
9cchhxKnhDvNoECFe/2Ya4/daSCpg+j95G4eFyGDihB0UOiGFDfA3HMIIAFpsb38
Un9jNgeNpcOL5X61vsbqe0BFnQKU1Uij1mfYtYEnImfkI19DqaeXU00PY6miab3C
mFIzEWsxwWwx18gYluqG43PvpXk+JpyiRIg6Axpv/ViUvOMPeiHz4kFqFpgVWyhR
cGxYpfIclc+tMFOSlcosSF3G/B7bnOqL+1+vtxpR2NoOGVkanPzMXLvoBoZHDwSB
x4w1z3QBL7IGSOikhAw202Tpef1z/NkS2BZ4me+XDycbu0P+plCltqTkqAxKYA4c
OZjYlngtta1wt5IsxYtS/bh/hvCrqHTsTuSIDR62btq6RKs80rTVvzq/GBy+rGdi
6ygPrjTTi+v3m29rk+IdwUoS0pE1hTGNlxQTOUBu0NXY4R1jIsxhW9n03d4pou7r
suUEqm7CkBAXRzMs3RINzkERo+CRRdNxpu1rm+7uJcTNJSQ146+P+FObwjRkHSQt
Fh1Ljm96JDhaESmQecXQNKLrbR7F1VJ7xTIrS9A1Wv+zOnnDRQSjdtN8ditZVk/7
LSriOYi0VrDAcg+thSAM+LGMBK7sGXrN+fKoWY7TxWs7t1/O6Nd9B8aJDx7AN8oT
PAV7fwpbGSf97sgPUS2YUXCWyQbn19+GrcFev70P83htCrNENy0NoCCpO216KvMk
Iv7w6U9wsXu3lAYcoSBaxr9KswOjUEX4T4TXgQniJfamF9GBkBkjtaLhoIoEJBeu
SuW0V/lnC2hcPo8Bkj+9RpkN1S02y00gyRJpUntZhhN5R+88QxuBFpxkf79OrUNu
mAdo5N45HGhPiCZEZIkZgIUPLDTmLvP72a32rBIDL+CuWgJOoBFI2HuV3tzMUSD7
BjGQhLySnoA28AX6BdQu/1+RqHeRJ5TejQMwNXa87Vx+irsVEPcT9Z6FsybbFWmy
MJN3KYRSTI3d1WSol1CLfCl8FnYQnXsVcjTrZrGkmQE+drpIoCVzfgfGM7mSoyUs
0AQldP92MDMHDsKEu94yuBrBr0/mVQmRtaDFerlkb0nuvkC6c9n22Y4GTAUjjsf/
pgJbI3efCa7SBsBq5Qzo/tss5t9ShRF9W2XOJgt9pAol+OBJrT0uTbHNDWvBFKi1
whvghgk2Mlm0NsgaVG5q6af1YbS2ninUsxLKDf9lksmPPnwEA/bw2UNXVhQzef/s
dIGNohaXEp2w4X72Q4PuxEJcwwt7hHug1DwbNZAI1ZmKrmU7cYVWtehjwG0XSKso
w9/vxyHhlhsrm/T/+Xz+inhloj3SHC7mM0hwhUe1ivDW0rFtwGnCyKEyPfwWik7u
cLDsKlR3GP1pIYDZAI7ZWMcoadsyKNF9ixmn775KiNcdR9xizfoky5Jv3kXuGHK5
AM9Q21FH99wEhukhglNn/3+9GWSUKjJdFtw9kWAskqJz3nKPEZapgkfyyYGB16G2
xiIAietwRC/rsBJeDxIJlTpMM0lDktgXxeH2SacdRGCPLBZzZBb+urXS+01g0o9S
qiFBj2jrxJa2OAxxx3dpDJ4I/HMud7yX0h1QZE00dA3YxDPLF3zzY8CYMI7PSHuV
w1WTtM/M9BPWlE9EWFwFwROFGrdXoJpdPHhyUBvUdvrnv7PTbUCHjRxEGTV7RuIj
Vt+9bTIBCin70vZO+/w/7G8J64coP5R4oQbHB+QIgBobfYo9BJHUsBVHc+XFvtP2
Vfsino3nfJQ+jJFdxXA08lhDlHKXliACBQTjSE5JSzgPvXmoliHQsmJGMEUXlPQS
pDcxe6vfwiDBXMKEndsm4yEf21ZMPVnBpstpV9HaFY20FxS9iCS7vuLIVa3YQ70h
FpehbLqcaTFgrqyS1dxD/3X/+1A0kJ+1FaxVMTJc9EsyWK/t4e7/ztbvwNZ4bN7R
y+kbLolxY568k96ndtwV5wIAVZS1XYy7den2pxAkkj38zpQHG1cpHaTdFFNrK+MB
dvfm0aANqt1ukublbOv8Kb6Dyyq4ppKYYugZl/q+StBoWPjTGYwS3TGtS3e8uqDx
SG1ixM+t7MvbR/4UwecspZxyDL6p9O40wRziyCC3Us3P8rqhBNg+FufUe/PGc7+e
jqi91ywxfef66h5rCtS3kqPpXTjhE8N81q5R+UHNUtZkjha0sxpHNcd0AFw5kDeO
CiF+Z+AzL72S25dm+XmKLXd2SvlhwpAZ1qCzzCMZfR6GynSZFWkwyJKsF4gY4HWt
FYnwDa2usgqzwCQispXro33m6w/46mL85GusKo6L/ieCkhOnDGVvYospDhBEL67Z
LKV8dti0b+24OuSn0hjZzzI4djEzgrHxEe0KeNaJf41MoMArlnn6QNkuO8MCDWUd
NshFTD7inY/avC51HrJxeDj+hm+3O3USFtppOG5t7PsUxkl/p1b/m3RhwIxc6fnC
tnmgZMrbWCyWfkCTk4wd0w96R/7fFIAF/6pXoUsb9sd76REuhCI+02CWrnljm9yd
R34Bax9J7EcszurjMdFnaZwmA3kI0pWtzPs2YWdNANVkY07SNvmM1ZwAYNUqgg4p
EGveTSwMX4PlDdw/4XZMsqlI4/QpBf9NG1VtALT96K8wS1xQsgC5R/Flo0UssGCl
4J9Zo4bEmRNfXheaK3Sj8t3dOYkO2qF/ApS/onOyFxWI/+4C2T2TG7+cW7ccZf/x
XUJsMzCyhy7oxD94Rzjsg5dWPCe7BAX4CwV8tWAhSaXuVs1UCjFWUtlu4AkaW5Lz
P46AHHMV6WrlmOsNcxzzbF8gZH7/F9vnLfoBsrjXnqDORVaQPXJ/8amvJi+ty8ca
tFXgHrQWfAvPb9K3o94J7HgGd6J9ghdfXOoSibEB36fFHcqk6qaUKfS59BpAdKm9
DKCFJYEdIEjvGsjPcKpyVzPml/f2koLMjzXaSoFqnME7tcGB6DmZeyckPIHiYDH1
tk0aCg65jLxpA+sB/uc2oIiV449zx7heevlMmyXxXqnhO67LRolHWy5PSygHjg0q
zT9PTLC9EpPstYsQi6xazDekfuq44O+l87bUu7JEzEamG0wxHGlTVOeLXD0hUJL3
hc0VOuTHKyrVyiBP/Y+ApOSRBMX/Lly8YBqfM1QcUQyYVAu4t1T3IXh87H4umk3O
nAvdh0fcf7OqfAK7c69q9k2Zx1R8Z1BAKSCWcPMyEz2tnRMweD5Aeq/OEDRyGGGa
H2ghG9A6MaQmsbqSHChFVciSXltOWigkp7JN+voTkPRZN5pMuuPd2Lb2mkmTsnyJ
vXp6nJVqScIHmkU2ikO1/4UDjxrKKDd0Tsv/M1FPNZvCX7BSjBlxQi+J7399voJX
IoyW8xdRZf5ZD7T8aeZKoeRRmX86m31oWj791YgZGFAVS2j1lqdEUNv0awtjNSxp
QkQmfZV2D/TOG9W9m/U+nfq9qBazneLPxpTfDMuUxzlk5pt+xicKYp91NWjO75eu
w92TXVVc4YyGylZIENu721Yvsl+FfZRffmVP/NnKCEsFaBb3rctuURu4UnZ+uJLH
MyXeOpyiRTNqEjqjo/OprPOoJGICC8LEjswdDGNytC8ZGL2//VHVXAeblyEMiS8Z
G5ELtX0kmiMvdgmpM6akNu5HpyyFkLQSUjDajRXbai6HXpQ2lE1RWivezWR3aLUa
htR8SKDk9Jm/gJLQyvuO6eOoG0o2ltWAb/VfFg07q8PP6T0ObeHQB/AVH6Tm2ivH
HU2uPktB2NF125I6T1APaZx+yg7kWTVEvzasL5C25+6OsqCe/AjjG4rs23OJFdnW
MZT86dIxf6Waj8xmPqHQ92DsEyxuI1LmzTDADqAMHMaOoNfOXOFXe7iDNoKkIaTo
7QdI3U2zlxh2Y4Yzk0H9nqETAgkMzM2fjXHpJk4rtBPf4JqZdFnzx9LHJIQJnRiP
RsAYIwEGYD4pe8A9RWYR+5WgAW6OgOI1ylWlE0m1RwE755Det2rzrnE/+fh43eyL
H3/V9VC2ygNFv97Wc5eE3k16GDYamCcqjnSMzqVEOvAXYvI4Y+EvdFUeM7d7PONw
OUMpQYoXn7+7/TJSGJib3SRyQ2ax6xHnU8ZiN/n45rmIoyjPY2UTZ8pbR6Sk+QSn
GcSu0f/JZCMRPA5yKScOGk1BroKk5dId4hg6hweuCGkVdhvdbpZC/NAPeTf16zRh
ygiZZ2550lAzdyiVxVqvr4de3StJaxbb47LIvPSh51iEw7z+cHmIFaNY16+IVpwQ
+QiAsmKdoGUHjU0itLyLxkWpLOn05G5uGjB8yCdPLDPKuGtPWtnPFjikG7FF17NI
xBod3H7byLsg93EW8NRcpH+cjuzmpkvXnHQQ9SrvTjknO3JIvXUuCAE/6pLNSxzW
D6xk7UAhDOr+bv0TZkAgHGNXyEMuIHx5P9vfPnPSGG0vW8JQ0VX8+SBlUMx/PoJW
nM8E4/Jyuah564yfw4KJMX0xeoH9VQU67NARnhQc9oxxWnmecwkdyM48TxT/hQoW
CRSY9LoXkuNlis92wlqZLDKc+XSvU9wcylWrSOvJza/yymeuI8eJ3usavSDzm42n
LbTv16XzJSSgcc+W4VmjJpEAla0kJzyBRNoV6IE0C23LuLl7zxPEovuMyZIvMNo3
y2ahMUqg65J9MkvpV8AKFHw+gcAdUa27dtd1LhZ4FQpPXKyXb+Uv7OJx6JK6uepr
qmQMzc3FAw3h1DW5Q5VNvKve8K8jkoqB0X8xLYtLsbzjbBvzBbCdQGyJGSuMOK8p
aq1IDJyknW0nkWWzqBHOMNYPFjk0ynm24/2kHMf9QAuS5Fv2qMISy4Pqqhj09cj3
3UnGlByUIagcM6z13m7B9SIcE6is2v5nCvsj/rkFZsiIySlQB768RnHRg62AFdGA
7Jtfgj78PPleOZVMQZ5QGjXkGEFQzZDJcfNMoNXHcEwxdJunaRXQ2NDU+ToChrZs
KBDlRtmMAH3YYOOdwobR65QsEvShrbGdL6SDTuwC1greRq56sxNL5LuatJARauob
cUfjmfDEmoWA+J0gN9dUz9jKAZ1C58LgcMHmPOoFp89Vf4sPLLhz3NFQLAS7iCWG
WyPRGWUy0AkI7DIk45pWHMNeLMJYKcCp17FyEfJcR+inEAvw/OnryWAQ3/6JQvxC
QCFcblMGANwxkoJmCSqD9EbzvsurtwDAEJGBSNVy6KgVdO36++oavh5AvHbiBo0Q
f+4h8qP/xq3AmBkRpm8scaiUPRIqVY2zRc2F0z78wIJF1RjaIqrqUL+0cQ+02tT0
g5Fsp/1yyd9IhvpcWlAv1eM0ueEY43ctX1zISZ1GhOZ1eMqsNeR0joxmdDmRKc1Q
chTYazh+0Bd1E1dNygHt3+bSxhj1Zbjs+Z+Da0IPdQLd7ckNxNZ7QIaELBERBmow
KJC0KpqDGbUPyKQ+lIHjFZkGSOkDpJ1zVMAYzwFiCJmGOqKdwACsUcZoHvRnrQSy
JI4Tfja8KPjyDjbJL2/V+tPD1OFEyX8OcvrpZbMobT8gb81MXCRKF80P+Ml2LTHP
ENErOfzGUE/PXvVk6YGgSPF7wpWp6R+T+3y3fq4JNMakKIFJb75V30oiu7XmZxzX
a/rZfLcQumtr6F/m9wvj1Qw+LFAga1Z7UbwDlfP4da5KYvkimDPHp8XmoqUXQbuW
NkEPJ/pcHHPvhj2sC9NRoq21gXlvdAY8a5nOVoN5va6HLbVeMRgp38KgVfS7ZIBz
QOnaNCfgU5Ts2+uY+RaD74937zUsnEKk9JnZyzQRHcqdDZQGEMP3FFtxINrCICh8
9x6ap1s9nhjstefSvdRIys9qIzGSUyBw42nEdO2W2IGSORrgkiIsxDOpiLz6LwwK
sGNWO4oRqkm6NzbZE3rEt5FW3g3hW/kDoZWnlkZDsbsEe/jBEelx+q1ad12i9XU7
EASXPSHIYCmWfJMeho6e9WgXcNJstzDzuCzQAJSND33BG/nFt6+UTfkVuU5xxp61
kq3FdArAEuP1As+4afRsxaiXBBIpnc0NJMl6poz+htGJIl/Lp2phiW2uPTwKG/Di
52o1Gu/jjIt8tljU7r8BrF9AAMy4DrBTJL8u7Fj36VLrQdtbAGh65zp+gHKaIiLK
B1QwSEtdaG9g0ZxucAuIWIYtKJjpyEGgWXxJSI0TUx19h3/gxAfz4TaMsFNNm1wd
yKFV4PbTa8r1DS/22E9vWS42BH5AY7juN8zRvi6+L58PtUKXqc0IPecAfjz08qfU
e+XUuU4mCxLdl3Rxm5K9D+TzK0+BntfLCVWyZ+Y7ZutbvJ2ycQWyKWJoZNkUQzfQ
bOZWdmhAo/MDyPKJYLd3xDCVXt78qawri3bhiTfzpTD8+MKshadMCdA8DeDhGKHV
Axib9mmqA+ruzia7hrQh6IZkD5smWEKpVTKtEMjvFJQYZg9Jv/qtshV6LToVvXo4
rxvnjSrqfLrmGrqmJVZWxceHsSAilGQ443uxo8kLcUo1irPLp4NctC8J5l04vLJ2
+YLJE1QZcXxKYj3Lo6BJAjaWcZKBC6Ut/u2b+mjTYXwab9rwjXya20iA/TiQvt/X
V3ZzZ/f5AZjZxJUV2HXweHnx5a1selzhlT/Y4QDqfvcoKkxdXMwP4+JHG28E52O5
7dR3NLocPhcR70jv/cYFKVzCVvh9gyq0NngWKwEpNODc4/evPhFmjCQorDizkgRZ
nxUkO54xntNjzCpREOFZrybwsjhL/vyO5vOfQOCvVMfk8XfIuAlRa4I3Pjbc49MW
L+YBKlMuAuI17+PH5hcIlp1ljp1zRwYgXaQPie09yHPngLL6fYQSRr14q0hqVTb2
C+UXRef7UskbphAX6v9yj6nkICOyi0B7fmTgIJmf+W8z+tRzKPPK+K5ASExPUPYO
g6UqOZ9vcLCrhiCPQtET/KDbzUkkXuTOQxkdhfmNIDt2I2LAMxZMg7aj1WvLL+IH
AKnqonUwk4Fco8pJlgG9htN+3kHtSbW86ViBN4ctiFqPn5DSNXx+75GZR8QCA389
ELwYSDNyb8gd5OWVcjbmu3Uyb3pbpzoYY9N+yZ3/Pt/0vx5ncgpl36OWNfLCf1xc
Uf/gulaOEk9of2nkziHQ82H4jS7VGiYfePMbqrI7r6wlQIiyP8B+BboE/2AxAXeD
ega/Mvvm/WOsbSm1NmtYGPT1OPGK+Lx43JvE4CjNE5gNMKWR3vDvRZI4Zs6VMD7V
QnqZdiWsJSom313GBF9K8kzKdg/7wu5gurZh7pmgCH0l29N9MfXd0stx7TAmtQ+q
5fBVIbxcA5YuANa2q9QaY9Se5SotblnJshIbwioswyGq+7VsAf8yCCzouZpTXonO
ugA+zx8efIE0Zz2NUXsh0RxRiTDkJj3WkToZKPJS+Gw1DxjxXfR5LBPOYxRxEpCB
8WKt0QCZ7WAUkd8nRaG/quKJomAl6+R7qKPipmP/NzeSG8WuKmP72umrMV9M3juB
G6GAzWiVLxULIGNcg++vxO/RzRqeDbDMetd4h7Wu0Dmdzj16s0gue5lamZsmCMD/
2tnbsswUtylyEeV54vBzLt4MjeRNbmbfl68WWAgASf5CTXfejTiDFmwagTLWF9iK
bTDaIBjf4MAxHk0mcvaDsx4DgqOP+BD89F5Nzl2jUmbB7Pp6cPNXBrwJGCBHVr5s
52wCpJZT4qeDuhkxVhPQe1Om9qPdX/ibVBgoKv5AIDTXD62Djg4kWk9IG4VNF+Iv
+3T934ruGtqws8F/hHq42ZaR81Fi124dgsJaGRQvv0Y135sxQP0KPg5o+IPz7nPs
HqbLk7wWiQk6OOEanI7LKwpmg4x6XB2+Zn8GXVrzh0W8iJsCPo43+e3whQp13gkr
FSWTl/NiiNc+ke5h84ozrsC5aLkHNW4m8AuySWfgY0ul89iz2JerZOn2t5GoNDI2
J/HZKTvR3Q14WU0lEjwEJKnXbVXe6uOA2zoszoPM4MKFPrs3G0PYFwJH1gsWr0Tr
orbM0bCf4VD7LXay6Dy8b4XLw8jKdaPyQs6dju1RDXbmiWAdPocmiBzT3Q/OIiMs
BHZWWo+0wSJconIsG6yPD9P7CRl6hzvXr4fCw7915FXaYPeT3yy/EnX73OvKnemN
vNqWf6+vIP8G/kk3iGsokEG5qNfMbnd8UXZTzLvvdZslcCJElyLG8Q05tRqcRk/r
fm7A8G8uPn5o4ebHP0N36SSXnlbc57nuGzppWFVwH6t3xZ/Y7X6poZyMovlaG/J8
xBQv8Useiyd+1o43m7XkPe9AA4pExJAKbZuzRKjgoQFUYauUlZvwoiiCuN1Hba/v
EBcffh33uEbvdn0fEQHcfQQJeLMDfLn8uCnB4ttRHeLLpnLhyUN5DSsOxH+0XKIF
3mZq4j6oKyOmfhASVefs8EbD5dXHYTAa3YiyN5x+Ha4GOKIL+B9fxYL5zHjbihKi
pp7q0z5S/4MOEPjN3xVZ4gS56TYxbJyZzyjImH1/v9R7MlFGo/a779eGgPVXn4IL
IRDTZibNxxAHPYFwXNOJBLpa4ZTJmwI/eEL2KHDfZOUjKQPJ+6dW4PMLNLUI3D3i
/EALmLHTXdW4rpqXMigXvbkR7kFFgeBDv4S7K1f0kk/g663cfGbSElcnhiQ1022/
bFS/ujLsDBwxL2SXntuILM3ycyeEAPQwv+d2r35GohJu1HsGMTyrqVHRxmVCX8Km
k2LOBbKuXUm2fqDOI8aaat0qMe1XGDgwS2ZkczRTJtm8j/eYg8pkeBXZCxyDGsz6
peQ55NyxSGZczcnydlA8JS40qF/nAiQneLKymQzga4phhOE69UTJ0JRfPQeg2QqZ
g9tS4hU5u5z/vaxjKqAErSRPCsdZ9DVubExGdIA0jjNtSo593joDpeGvLM4DQczU
CGkgFZr0WlOKZbKoP+FfPBkwqD5pBFF5NPrpqBtPthDfziE887b1Bqudmn+KfjAL
NGMwKTRUs5NDvY38GvJ93yc8RlrOcGmZ5JdxsN1/tBgTMisBGO6u8N++Fqyd1CVR
92/kUv3b0yrnbmfVuVD9E+JKiJODb6G3ZZx7DY+So819Xm5M1QHTzKnkEDyfBr5a
x5Bl3qg9ZUU77JZ5ns6FhC7ePLbF/bHNFQF61oeWXlsgZVGHvXbitvmXjANg4LvH
WOzNeLHbwWO/vdLwDSVaAl0VqapOBCsmw80jVla2fca6L4TMDOMhYX8KTLTYy06b
7kiKKHF+E1hBGFZcT+5j8RF5u+qsxCClLlWvry1tQNo+s1YnFR666xA/ogWdvQhu
ao3kSNPoJbtm8aNgLbwwFF/bT/uzyZnhvaQ9ly9e4Ldci/AdzsdEJC0KPMVRDzFp
KSkNB9eQkOKjUpFR/RTq8NiS2lcZ37CPH6repDdcDUJzTNibY7Fojf06DtdhHZmO
c1nD+wA+6hl1G0/u1kFjbpfjlCOKBqfUM8VGBUvjKzLBAP+WQK6V0s8SnVdVgeKH
jupbsp8vddUtRCXZxh+Ow8cDOzZB85HtYDvy57OkZFCishImnqac07jtLnGlCmhS
ytxdFIv3mnpJR/HuxqxhiD7+GY/maxei5R84ywqwANFkpxu1z+8V6Kn/kiIqkf7I
edtzXyQs3USjqXgbYTTckDmPSmFwxzXITPZkcB6tVbxSlO9PS3+2VongEDCxxQ3X
arrMwayiwIghIRV++QE3ucccyo7H1bhzMhEJefOxleHhew2MkvexrMQHNKBchPEj
6OfC8V0X2QwyFTFCRIZU8zhaLjezH5eWT+ttR26Q6hWmv/wxEdF3OIGB09eXa8B8
L1s4trXmVTFY2xe4tJ3S5GKORKidyPJwH5DfGvSZJA0EkpE7+tnYCfVj8vP+BKAb
GSq87BijP16NPAkHA+H5r57AJx1nrVQun/dAmyJZy6E7lOm+ctO19d+erw6QVdKn
VuGBbD+NX0JxAbKrL/cQbfucPQLrCt8Zv76BEpQUxdwtNb6TcV4Hvdur2RsJZcxt
1Bct1pL0hbqJT1pHrzUWrlJyvbO1gSYqZZS7Qc/dGuqN7ki5xhIV8Mg+8v8eJifX
X4A2/5ZZefccN6fX5fXMkJJjmeKmnGjXvqmtCkXIbT6/tu8zGzmgnVj+d6IKyvr3
vAu0I3ZIYULy93xLzHAUyzxCPyTXU1+k9QUIVWrbFCyIChLKHMkRyLr6JIP1ZoyG
R88rt8e2p17argV+FxhPM++4DwR0HmZelm0rPL4GdSoDGCsODDmZFeh/XpqdJiaC
v1M/PV5kDSUe7IFInPUMYYF0YvLnNZJQe0uqUoV0sSDKM3aXs/1smEnLtOd/OOSX
qaBuoT5QgbN57SN/01z4sWo0Jtym9cgrfzm7FeJ0smVdEb5JnYQ2jcr/es+zEOqZ
/XytrWHePwiY1/FezSU9nPBThLOtkAV6T3ZPFJ6ZvFrHqBh3RX+q1Sx3HeAlQ+l4
729QGpa7Eo+Ckk7d1SgUkfXklJE2VS4LuKtW3dl6pvNSzxaondBYHFaTrHZ3JZ0d
q1lQ8iXs6N+sUWD//lZtlWDSM9YmBG4mm49T6MZHDjq+KbhyWo/NiiuBRx0bGvGb
xy5EZukZ8C9qjaZytzeO4p8SQYAkx9CrIZ2zTM79EqaLiv+mvafUY+Zx1f12R7QO
0WEy32YYdHj6heOPTHE/m1XFG1g7mXRzPeNbtk/D80E0g6Z+do1fo1epsuIRJxGJ
tvFFRGIb4bQxlK9NXuPx3klSJF0Jw5VR0E5ak88bOP3SZbc5hOx4/SSStE5BQZYV
g4pTScHzJOadyuCIvL3oECqttWY1fkQtmAQUf+4PfT5m0BPkSDcyDJpOIgLw0U0p
0uNbJgNkVNn2WLx0DCsVNmlmtKbMngUY1ea8fJ9Ok8bQ2aVOipPptKfpZClwJa8M
AoDyDT/h3kMwFr4MEOau+7lqkJyYBAzCJeGyrz2FBhPjhn6pIpXvIJlLV+5Iqy52
U03GIbvlrK7F0sOyNn4wnXBlT5hLDrFc3HfooHadqNNyrex2GuJx2LitpH59Glmj
KlXePBkyl2bnevOIYQ/kr9lk7qbhNJKCeCBIteRZDsrrhAJ/4d3YzWvH7lOBQE84
jdn1tzTTa5MuNbHlp607ne/QZhzFcw8YrnYB7MQqJLbSWPepGYzXfvxO6x52wg9Z
v1Qgb5jjQClhkhJqNpqBk1W1dElKZJ8TRXtZMJZDdjQ12Ip8bk62MAuACSI3XSkS
Xqoj7/A5axlAO/4L5BDs3I1mB4cYRyLoiTArmFv1/NzZScHw018o0w0uG8VOaMpo
NjRmbEje8s8DuCLETg0e3qB42fgN55qfW2yq1fwCRaXJBXBXE+CtXMwiMk7iL8KQ
/k4lt4OUri8tabh4I3xfoYkIdMZnmV0vmJ6GZW/LiBdK7CVO8pUAPeDl/MsRXEje
Vym67rwYEymvfNk0XGvpxBt0DqPQV/0iqOjnwBznMVTyBs/RsLKaFLKIGqyA+53G
4sJCX8YNQEbrXPJ4JvbB+FLF+vRhy4ZUENlmYjDBVWhBhV3vUnwy5mhmqUg7rwXY
ZFN9pSAxHvzpIccbmfj3Cq5SXMcbzUHJrpRpn4c60++V8/RlfRhMo2VSBlmzvoHo
tZTkt0BjtIoYiMH4QvX2I5bzjYc/djLY3+V08CIlKhSyE2jIa7dY0kZh+WnqIp76
UBWNCamZaZ9LOqd2lCdzMDLLOzEDDlYfwNhESLBsUw/gRkKOZ313S8SDC+0q1K0m
GG9V8XeyPCTZ5mkPMhSFkN1GZqJOPtzbdRBL4Vt7E3x5Uc90MP49Q7wJecYRvRbx
+dHMmq5DZyJKX9jL2AzsJqVrBarV6Kus5lz3pgSBEENq3fdzLUWyDDzRblLAzR1+
RY2dn7Hco2gD+5jOLTu58nd8w3PoVNO6eJ+hArvKXGpubJXztFdXsaNuLM5jfGC/
xlcMx/X2mHjQVXd//ttMwZmNSdDmkrbhwkYRouzXO2HfA6FHM+l6NABl24p+tmiZ
vkKtW7eMcVO3NXSpwPFrAYY6OJgAIm5fyZWzhjsuwNJUSaqoXeCnJjb6DvmQuMfJ
74yK/gdCZ1ui7PkpSBUWFdvQjGr2KdBJzcsfoqe4W3BN3BIIzNzcwP2lJlaANV2f
gN9c6XXlB7D+kA8jIleCeEvxNE6pdee+M0qJLcdDaffce4UuN7FEG7tmCK2qe9lB
/7YfL0BhtQppkwlm+kOXzLVWVW6Li2PYgL+ULBN2vpEhdPQDnzifuGbKHGpSct71
4i+HBFkAsv9juXoHBiUxLRDFRTfnU92B3kvG2rX468hhqd+Z5M5HEPlPCRUrY+mO
CgLAIj+PQdUuG/MJ16gwTTYRAOwKKErktzrpN2j0magle6YcctfdicKPv6dCG8o5
H5w/+iPZCSZhBAOcQJ1gqFoh0g7v7+CORIHm1goPHl8nXQ/U0r73gWqc1VxuU8PL
NeaMkD2oPKU0vh5PGosz7Ja0Te8KB9EkZ/SWSTI3jQlh7x2IHrGgmJJPdHGsEm4y
DDwJ67BsssjLjo7ZjprKh8LovCUwXqv3nVTgTp3/YHy6DoN+XVL3dhgT79uV1OdI
NdXb/aL3gLtLD9hQZBQfa3fkL2h772vdXX0iDk3Tq49e8hVjahvH4/b8ZYeJgOwX
YdokIE92jCb6hmkt4pjoCUhN47uZU/xi2+Xx+EIWGN9Dr8U9nSsaOH6yh1XiDsym
YEbY+4bEuI09VQSij2UTGqnX9CO1aWrDvlcxG95f72JbpBmbrHX8p8M/JiAsS1xr
vDLnxsfMJGk6aiU8E10VrU1bbuW8smnFPSsRfvsOPvdvPRNmdXDGpicqT/ewoF0i
fFbN3kTY79nF8Qzdz2Dn5ACJ5XfSW3bn/c2M/xVOfVNvCtciVbQw6ansdbKoEBHA
sWu8feGqohoMj91OwP6YfC5O4FKUFamMLmyueRpUc6fB5GZNmNuQgSTIG4Mr8e6Y
DWr+5392alSR0NbMhqg7uzPNENZZk4/5LOTuNo0R8goMaZT7bz0iF+1LrHihGTMK
3gQ2Ty9fh1LPBsRp+0/QkogDM5ePJGPhMo34ZxUv1O+9uTlkPOqrhy1cT3NYWGPY
abjBy/JEwL1pLPm4aqjAHcbExNk5QsH4GwBdxLYZ9Hy1+bi5pUsFSg0mmYXk+TF0
79ATBBS10VfWBIslRWUUG6XONFFJ/hGwz0XGjhBxd8E6SeD52eo9Y4bjU3LxR/e+
LDJfRz12Xrf2cWkayg9ZHchlMYpAxPHI1m9o6aKOHex+vVCqe2MTj6+OHD5LhMRE
5MfTOeVF3LF7wxPq5cQkJ4aPsQ7/uBjaT1yZqonLfAj9fKr0fi9UcbvxGOFOmfNp
WCl8HEuxj5UfCkHJs6I4TVZeaiczFaU0aWJbDusO0LQNOL/nvu4Y63H56eK+AZNs
85Ro/hKSDE2zJz99SXihdKSnFqCfIaRk6eeMrfJIhoSnikLWO29S/eWJw8eHW4Ty
AfVuRFFQpOhQG968hsPx0Qa/z3/ipTniVCw66pUdB0bpUitaB3LoJvnzLW5oacVa
0byjoNjIJFpnFcG67kOdFYizAkAnBFlmp+eHKrK04FBl2/ML35cKvA+jGQ1S+Axt
cje+V5dLZYaZZ6Fij99AAxGI3dA0XKemE0z1eq9WwPNYQzvYy7PIVUL2EGyNjBWZ
8U/PrxRiL193DTzaj94N89nDvoutmGQohRVlt8c/VjUg2wcK/uTB/BRjHTYshqQ0
CEWoSYvKJtw/RMLtsR/ieiCIAnwuw6INiLIrCfku2TwSlA/o6dJQocDFjmxVLTPQ
1o9IktQkStvzsSKEKMS85lF1HrE+wLMMStUpN3ZRyMkVUgBUGLjDrk7ymjY4Gd5d
K4GXGqr1ojFaQXIGhY8PpDC3kSDLqzsex/qD09aMPHDVMP6nN7RPeY1p88stg1MC
3zVv7DQOlVPszKYJc7YmMrNAH6XpZuOklNYC5qItzaKTGJIelUQSQNIE5SpGMym0
O0Jr2YrMpBpWcjp/efQF+DiH3qChRYJM+I6/JhleuuipipFPVTc3YiBadjs3NvZS
/rrBPta63W/98vXo+d5mgY7BFq6qKPf36RL71t0Mc2NcPkZQODCMLtazD0NlL//B
CHIxMl7Tbhnk/AeB1ribw/oL5VKOJUpSez5EqgRhA288bhQ1qa/Kb7adjxW9xwlu
/DhuTECSdQVwJstr7hajeOSfoada6tEvBwSl+IhQASvrrS0hpN3I04/jgMb8cbxM
WqyxzWMq1RTWoKEV9w501ZJ4SrXiaErzuZ7FJvWULYh6V2jHWjmkKU1HQQAfFNkq
VujA9bWTdTZcZiudSbv2pHBDa00a9X/2Vfz9acRTTNGL5zWlK2zNTueFVCNmKHwN
mQUXCn1XPBIzwnLjVVw7vyjnID5K+4p/P/yskzv823KVHXvuVrh9j9qaBkp8zxVK
ceT6vPNvSdMJ6UteRAgGmsxy2SQJVYY30d6kyF55fkzaS7NhNnlRmHFcDLW17L5E
k0Fs3Q84pAYAvaR51auJC/ykFwRrwWZ/VFgTrQcRJFoJ+La2f51CpzZriSVkhzTu
P1IZkeZ9uAvloyVryblF2R1NcQ8SPBm1Q18nUhx0wq4ueKF7jqjRLIHeWmZeNziE
Td1IZR83xKCwhUCjNvy2c0ppAuOtPC3oZhdHVJhPRV2knHqqgrkLOEYyd6do9oKA
JQIIHacKQySi2JEEmea7j1neKnl7j30ppNFViccVF3yFErj6WK/9aAJBbVl33f1/
Z9a/rtKoMNKPofitkwV5j1k8YWDqitYpLygkymOw97A2Luh2tP2HE3p6qMqIPO4Q
arkkifuPm0owdlKjxBGqQgeuVo4v2/SWBDJlXiUu/uFcNa3zl9XXWwzbN0XIrDt7
6Y3M97NofS3eCBL9hrs6OLe+8w2vxctSxW6varFiFzmQWKGxUvkBKi2NoihOiV9P
PnrOOpXAHYwqp9Yw1m82G1CG4fAA/Sk47HEk5VwpM+xw7PLjHT1TB/hnNoZopQHJ
qC7jdH6RlybOtq6a2QM+Bf2zS7qWCUU3VVGpU0B84XvBQckg1hoj43+7cvSu4HGX
3GdnMxFpK3xPV523l427sHufoUGxhJnCPBU4tS/m0XQWLqshBaE5BWiMSRp5LgCm
QOHUkAxnTKhlRmR0cRfJHYYFvy0EroFMdPiWDWUmi9gY+I0s9Tt5B0/5wv1KKO75
HeOmtEQj+asZdBkB1xCXD/bsd6yJTq9ma1kNa2X3SXglM6JX/ZPWyVhr1klAmx4W
YyclnheIHJfKqplckXnylBrx28E5/5ftnI9C1nfW5l4HoCCMR/icG5v26BGrvEn/
+7jvYdj0OdEoV0ylS83xE87V3xH/ZGNykYZWjkHq7pjhFsNVimc7T2KTi8SywHex
NluGUxRjBLwO8aHuXxa6cXawpbvtZ02CCeGJ9FiQBQIefhcj5f11QAOPff2PQPEg
/schsvnRkFq7ZA6jqfvQtLe+WyfNFNN4/F8Bzey+OQh0Tc3wR7AUjsh13tVXlL0D
AnEAPxgZHdrAvUjBi/reR5VYa+U6tlbMqBKacNyhR6cr/dErrH9nGirIiQTk3kvW
qmg5Xj6lQ7WcyqJhq+YymnhvQMfFzEJqMRgJdNMfx7wCr79spu3cwkSefDNviN7K
+sJh0YT7dqhj4hWsdiHHuSszmhJQQjgVb9rXJmMxrJMSDnHGTgAZqs/bcosmwc9e
VfxWygJfd3R+g0lq3algiSp956Z4XZ5DYkVc69GObDwHCoN4G9AxZW3cQVdiiUjK
ZmuPVjlNtuDvezdWoa5WlQWgVb5zA/Teh7DCGlttttBDNIo053pvwSoHkmkE1AFF
IH1gbHdyDBtvHSAxMVkd0d0or73KLNl/SqybUY3UnHcR4B/2yJdFjrmSZgJsvKPl
3FB9Yuvblw5/o9Bw/bWhbj3EPBru6xUcKXqdWAZBDVInmEytqBq0+zpscm6cdqj7
Q6BffP8G0FrO/4fo0JRtXTSSxCdp4Lj5+wHOUPCDbyKWK+GwTrCjwgP7hBKy68Za
FzpSRd4U2qTG7wPbNN9YQ30vdNbtnHzayhmZ6NrVeyrtl9+81a3HHoDZqB44IwVb
v7LnUAnoAJGjNIF80qO+BwGkrtZzb/VJo+gAIAr7GKJStoI21IQMOVdiPiqgoTiT
twRV6gFke4ZYb83jGi2i5FBN7LioO8mMjSkq1IIbrSrhoD2BIqEIzt605mgOWj3f
b/LotGRneiXDOtw99aYs8+OSTbcDFuuSMOja7Ccjh/ySi7hKWHTtmAUCxm4jQbiA
zGHskeQ/T51rRS6sRubXaHOEq2IMSIZV8dXplZMlWTNhzUV/KYzgz69I+fTspM8o
KbNmtiBy/Xd+JU/ByU0RnKEWAc7VFvLacDrZnwIbO8+ERkmgatChGmFeLyer8C10
LWoLhlKEYC7FP+Uh/JgvWsFVqWyOoDfxpXpKZ2iyAyBMsZ+rZmHB9c9ieeZ3YH68
U8l8rqEco8Zpmt5vdBzVEWKpnl7vHnWHaqOnmNZCNTmRMchc+X5Yd0LLnIuyp37M
aG+m7BEo4RuqyU2sjknjC8d08sOuP8R4FYhOGSWRSJhWY9WsjVy6/PRerCK97FtP
SFVAn9fdULF7lG00s3p9uOfLtXKeoi8Sv4XSiDn3UXVkoBgExviiEiU+5B7pbnlD
4D3k5izfj4WfF+S8kyLHXheedM9MeDkIVCi1mDgKrCOH23SQ2msqfYlJuuyMAGp1
2L6GJSzeBSikZCn7OJksDda4XbWTqYI2Ns8fdiP6ngZPZj7iJ/5gYDiTvse2SC+x
rR+bM775q01gUStsRcJbkyeoSJVrmpqVK6uNT+0DVK7E3MXAw0Cj5iNR71RBG1q/
EgS9g30dMug05MeLHeEAzjRpyaJhDJ/gHlKjKmt2LlAbA+D7/rnv4NTGCYhOB3yq
nDY8zKuyGJHKHVCG+1MMjo8GJRbmWEQ+SCq29Sz/ZppVwJY0FjLio5Fu+IJok8Wx
yY5IycB+bz7AXOPdr8fx0ao6vJgh5XlKE927KNteJ/cyvNy9RM91H85f3vg0fcmx
E0SKxXykFzM4dqOU108CXxOKuUITdXpIGUCTXJTsacbdr1eMQapxH/9HkJbQBQFD
sg78Btd9uJwLKO+4VrZWNTwW3brzEpuRpVgTLO1qOCYs/mi2juHBZ7m1uYWTtmYF
Dgla2iHwxrn+rxEpYuv9FRTZpt11JpYguLoPcApTXL1gyaHG/u6autw/Y1qiYfjs
Fmz4/oGlGpNCwad8vdOK/dZNak/MmlENXUVBKhVtLOFyudXlR4SkwYf5nHrXrAqS
HjAmBRxGHFBk0CRvnqkZC9Jb9iBRbB/0FaMTfyB9rwZsfgqmCjIfoqLzyLldOthl
3s9vNtcDRyQx/0l5V4OBCkDTRo9zQcXlJkjbfsUdgnTEztolojLNQWSGSd4yVh2K
qetKM5WMt6iPNZGhvs09ifmq6JmFBAiEQenrjSN9K08ioJNPUvzlLpqwYlcX6muw
A+4ExgI6sVWoK4vK+xwBwFzv5HMpHCcLyR6+4oI+S4Leg+ZaknyoOB1kGbe17gTQ
Ev1QUq56IMaUb950Y8fjLaA/5QOPz8sj5AMednrKoPre75FL7Q/nPPf9xqQIDR6M
tp+z5I8pCigUvRoWMGfYN3Cktyln6H0quaMgS1Qd6rHnVjAeclF2ghzgskGm15c8
JHP0KIPqG9tWtWDBdkJ5/dZpjgy2e7PoyJyoChA64HBXl03SzIRMMcy6w05s+Pl7
3paMEF8S6T8oCuYKgKHs4TlHoKR7pnD5U9UQVSvVqVInx8JVPl2dgxt3xYRR6ge1
OVONMFFOxGYyKGUfPFogBrNMLuZyN+Se8YnRR/zmHN596Ol4jT6/gG2efeW7ft5s
KBM1qsDs1Ce0GuutoKfkkEchV/mPBomOT4AtgsiIx72B59HQljkbRP9MQR2RmuHH
leDnRLOwzu9GrMTZoCfYJNCEkblj8DGRYTNd2Zm5Q5iUHydmYSTNmTmnVQPS3ekM
iL1jQu7UCTDqQxD3VlEobadaNvzU/96xWhH60eggzayn0jPaIX4MlWNHuvmsJXR5
WmNBd3wSk8Ga9iGHFasftPaePDsMEGQWIsrWZkpCfa/Qaf/NaE+kvqded3qoAy6i
33GQgiL8IfXM+QXfIhyDadu/RgjQJEJXEMVoV8N4NfKZD7zbIu0oS2swbgAsGRwE
OdDnoB73yYbxSwBsYd1HsCveTZPzwYmVVeqLYyjroMZhb0NAIhgdGTYWoZu6u64d
ABbYAvTMY954iwunW7IuCrh6lRa7RUI4Kvun+0P5PmvN33lRr7g0A/KNEUJdBLlQ
pYtlGd7KcmILH1hqNo7/aXUMbto9+DI3rTNTznOnWzknYX5/v//Mn8oigqZUkI+u
pRtEZHSHTjLdEU9TzVU6FSySGwcGmU3QFMXo/RpnBdKxcZz3wm2g4XErPJJvXpQy
RKkjB+bItI15uIV/rpCUGMPqt0Z1ObQ8mt/oCeLCnjKEAn5sLXvIT63t7BJZjpJg
2m/UVXoEFNCz1XhIYJS+ljEVcYKogIMqQo14bxQWcXYanQqe0Sq0nSxazb7jvyXe
UxvFBpAmPVxphfUHHpR8l+Ah3BySnAG9uu+3aHMIPj2jvCjRpnzwEpl1AYW/MY/Y
Xa6BoreTYc0E/t6581Q7faWMjNMe9auyLfYi67uLXYZ0jD6Uj8Q52CN7kQsHsV7w
mTfmzSG3vxMqGeFUjMz5J9dFqm5Nj29QRyCTNWIV8luzWjMpiZPdEndD7iHEpTYu
uDIEuOfYRx+vYQnGn/cYQznPGE3eNGimUYQoaQWsTXyEdjVym2tcGho0iboEh6PI
LhhwHmZJeXP6fkfAWNs4OFO8SXI65fZvZedjw5YFNvUIpN8k0Pxw27NXXPoUVSGa
CqvjGQzEph7/O6L0FAXRjopIY1vwCe6E3jyXhuC5uE2BYDxytD/DW+ZtJf2z8sFz
0gZX3zHMb7JlOZfWtx7BXIVBMc0MjELCkVYuh6Ferz7APgIBLUaJrxzbEhtFV93Z
MN/lYwqe1xEWt22JhCYgbehnWC9/IfhCfJgz53TwC2Vh+A2oM0aEK3U5Hef9+eYr
HRkcT+VK+s38oSDJgWT0tRFYG/bxsfmXCeWlkIA9ZTBbPmBheOg4qNTvtCvBrHE7
JODhWm13G0oltJJgCJTsVky6ehviwNWorFy1XNP4oLnuOfJkwrMsMAixOLil+u+8
OKcogSl2csWbPsNoA04bj4QZmYMsrpZcGHHjzwGGVd/XE77tLmd7adbML3wlroqW
/PX2HdQfy87eAaexTm3v+dr34FqEkm7lj045pcbSPjShlqzmupVcbpEA7teceZq5
6hk2UWZrZVNXgbLQI8/pmclYxb0AcADcjONTbwW3xIXzcfTzxc7fUhpfP57hdMiU
jNjiuVzt4LI5K5/co6LRiCVJpsn3TWRCSaDYzg0nZ+3VfMHp0SYlf7LBiIsEnRbD
t7Kl69adgHlxiY3Fl2TyVLgdsogwrkYY23kKhKo8TkN+nRNEEodJ3kXLHgxy8VOT
1APMr32DMfml5QWejmh4d7oy8BJPApgLyigXOO656NIBhRfGe+dCaWxvOznR0aAf
7TK/L1aJCW+/ut5zlNEm/zjeVm3fPlYXVTw+LnQ/pk4qHia7Z92tNyMffifFmWqE
s+RiKN3WZf1iUnyQXgXWvEBDoBCj250WP6IQQ6xRepM9bxZztGWvAr1GMxr8RAdD
zHJSmoQIKGoWq/23uhfhUBLfeuneceRp3o7BCKeUGHl2O7eZ3PkclNGJYE8gvVeS
8UpZyxuTg8JeAWNAf7m6IcIdJ8ac1P04May5kLpX0LWbCmWKfdhazQl0Mka7BglS
VWaylG4dY9nA5g7fKrDv09OmyV6orO7KfHNxcRhXxfcwyhC6vNSh3pKdCbYz4AXv
4Bjv0r7fndNXKBgsvPtO4j3zOT7oUOgBeiK8Dvw08/DubRf26upNp/MqNXN03F8o
sdWyJO/h4/VOVX/g3hK66yqbmQKgtRU1uhrkrrjStuRZhzCxD+WRa/Crc25CmI1W
/l4NnB6+FYv62MrR3N5LrN3Zp2ZOeTdYxd5m6zKDBxs/52gbX/M/kipI9Sp2hFVi
z0wzMOJ0mRmlU7DqKYEV46cJl60loY3gSTmu3ELgaT1bgJloQmV0ZaaLy8z8node
JumXrepd/pZ77COZKl1q805qfNVWkdZbTZYorP18BVQBX9lpeT4wfghh6bMyLhln
wdATsWihhHCUx9aFROiZPMhllDwuzx7ROVwNiZ3TRgR1p/7OJoFFKb69t6y1rnGX
AEPU/mg3guxcYdmO2/wreNyxQb7VuYvSRBYlvIyLtPL2QKLiZKwASLhZiwAhphGd
CXfL/wRs7mg55PnsPs7+SddWsfXEfIoMoajiEDimx/Rf6aJXhuTTWHr/yoHgP7iG
yHqBMww625+/S0dAIc+Mg3sMMEMkD2tZJ4Kf0xT6oHxLFh5drKTN+gzrSQcJlTYR
OBJifmSi7jrAEiWCIQh2Gebb0+M5DwbdiWPGCOZzjSUNOX8q6/KB9+70z8yNJzr/
cAmbXdKF+fjOvBma4AtKh9Od6NTCWa+1OrpFHQ9aZXkFh4hov9n8G0ZaK13nS2U9
WioL3RxkFKz7tspZnsy+g2rl+PWYVG/d//L6OgNB2WEl/63dbe1QsbX0yjrUqJjU
+4LS+MoQtC5BPsPl5wuVu6nPOTVfPLuDPXWPX078v7erNxs7sfnrrqEAxnMjqb8k
2qpWfiNcfoQFeg5hAS7CYhZFbTSR8py1QIhqmbjO0XWxHy33bzxKcidfv3mUsJOt
sxi+U5XK90rjN5hEPmuS5eXGj3bBnqiARp9qW+EH6LP36wnf97QgCSw9xaGUuwnA
5shffIhrd+sAUixaLCz1h5vULTW3RZmCEO23bgE3gbax/TN3Q7XG2djYU7FjiFQY
4saU3qEcLgerYZV5Uw0X2o27Z5wZAQGeQRgTPoydGce4ObkmcNozdBK/Z4xRutfC
dkdmPQ8p00JWwS/8yHvNSEIs8kyeAGJAvaW0P6axI/bHFHryGQdnoOdA3BceR8m2
FKjTARDkW+pu5KEupKT9TK02NQM+f+odvu/SD/WeVJbRA8kSdXvY84SIQ6rkOREr
lxz0oT4qNgwV+w24ChXJxE65X+f9W5dCOQjV83Q5rFXEd+MCRKZzk4vhsQ2T6p+v
OIB6OXTjouOBpBY+9Ij8nP442wi9uk51NUOx2jfIi2ShFdgYnIrSP3RKs/7twua7
i4l6GKA5MTgExGUNf6T7duARxrLngXQP3jeZwofMthf4yLdq5dXnjDoCJOgz5LB0
S8X8WUyAHXtFTPX/CXosXpDGGZTujz+392+uXGkNPTfSn2nxYGBwHR8dCrhuqYKI
xy37E7B588G8oIhpVi9OSkZrrMPUmRmDAI4cjeDLR88biomchsditVwF3AQsceJd
wPd/b3SXDq9ji+NgR7BG/XDg/2Hn0fHDXBoiL/mPsQ9JWFDojVFMX+fCKwcuI/vR
X3r66As3foE1OODv3xJgnkgkmPmn8phVXpZ5BZZT1kwN3LTusbH7UTpMWwh+UPWF
RdwVhVxcjepQSkAqvVosVS2DXSEmmSZJXW55jDA3Nz5KF5iBIPakSTvwrTf8CEDn
Xxibw1aOVS6m7/G149C27KuzKJLXk4a4/pjXj2nCmYhNpguSUOY/mqaSoPxGOLOx
BOehde4gWxNAhtrxcKg/A8VOGGwUKtmcTu9FBkddarIxMvQMek4/NVW52o5tAtlK
A+nfjFX0QsvoBrDlJ9O5xXF5uCAA1tvy78yKAeet20Fn2iYkg9hGZAzImc/iFQc1
QUjHZWwOELge3FkkZ7iHxKUI739gfsRd759MDbLCY0eRzVeNidTZWhvI9FaP5r1R
u0deFGTof16ffMLhafatKkAxtomRk3u1Vd+Mr7ew7YUhJjuSqlZ6jphLGZUeEDN9
0DhAz8UEde5Mrhcq3frnAdqYSBZqGATj+BEQE3eVt6Ip8uU8k52fAWh2pjhzjOGc
SSvkEOCKAtLEIjuha0seQA28V84ISoAJtYF6j9a8EfjEZvjuChAOtRf4jnwHs8c+
jR+gfytCMvujeD03g4Gpau7ImjrS+uk+MfBLea1mlQuYziM2fgPsl38pYKQvD4cf
/+5tQH+ayxcNhEY+Wjo0rQbz9uvEy9gGvLGg6uXwi2NV7PIWF8CiFx35huRYK63H
fZ+NMMDgxgckk2TqVJl6wUST34El+vO8dzJ9ujaOfqrI/S1Scb/8K6TbXEtVvF75
RYWzVL1+bLf/ZWXIz7xauiiedCoEfDyxyQcmrScfEzo9WtCqS40qZzGnVdcBzBxk
bGbPno4e5ocQ+kz4XfxZuEQjFtn0UuJhuRyAqcOFx1rwP7CeO0ickdPGm4kuRJF0
caNFimIHNiofdbE6bDo11vrNJXe2HaFKuyFrg0Iu69uu+kMz7BscfyrxBTJHSvG2
21sOz12C5J+bGHd14XF2U8zlmI+834SiRDhFKd1imMfGz/GXKA5FH8F+b9Y42tqW
Fa2ggp0fQF5+e/uHyi4Jv0HBTyibJYN52sVaCij8r60sEE4ee6vMWK7ymRjF4piZ
zRfNgk5qplpGz3oN4la1SXWf0EEkTYQ3wWLLpmZC0OUd9XrBw/1ekU9vR4YbEY6J
Wj4cgDEY0UopAh3PVu6dDIScPkvD42y2Vo7bzRlmYlx+1Tr4JA2ovkjJJPGi2Ly6
M0WgsSGC09nWMmZv7jua/3gCbS1CeZdi1t0F2K7/Y9dxCuHh0jxbO87admR1W1WT
zHPQhF0c7LUieePtUNFnDeWhruII6WYpra93jpoV3gqLdlEdEu2Dowwem2x6ECSi
1Fu0IvszAvTnwKnw/3aVnu1oRMf7JWiyddJgSpF3Ij5ibS2vu6jaXd4eMH++6NcR
fwDeN8pWsuX6KJ+jTB8yLRkk1vW/XacJCVIsi1furFoMO17m8kOI84mLcPTCBZng
Y7tWbRX+LYB1eQd7yAflK9PO8V8LR3md/+f83gbAlh3vIa02bViq+SQj0pblDG6V
KjeLNMTAK5qyN3HYzrGQm7gJNYvNXdmqfexHaOj4bZsq0M7vla0RyPhp4kQGgixt
QFYsHEWBcCVypOOK1lcVX+v9YFFSd7Fu+O9LH7IH7snzCzYJiMeheH3nv+l29hXl
ubfLZ9InA8fouQ+6vHKJlOeNyG8B7KI78swk3vpab1LCTcZSbcIhVegNk7xZcot3
dqya08cJYW5I52jNvJtMYCQU6hcxKQSJNVc3CT/jG6pJrcu9DTWrCw2zDLF0GEtg
hO1dRJ2jy/O3TiAa8n0az0+BWcY42O2Lzi0LjcYIQ3npvfMSiOb8uOEznxsYvaHF
WBCMxG8JDqQhMQ18mzQbpIRUjgkCSKrech2GTlxQYUFnn9kLzNGSrAoeWtBSSbMo
TkpGW0sJjbKYL0barpv47xIrk8JqIYQOQ7CsN27aCGzGp8MmjLFv5vT+DnrUq6Vk
ulZIoe3MP1HhdWq0JnRywoc0c8TwjtzYSvjCnpnqmnuHMD78WPBbZGZ0X0LgnCA5
pPouysYDt2wl+rIhg/mvBxLtdgFoZJ5GXH7/CVPN8+tNJQfXE8Dxk8SSpOXvMLDU
KH5LVBunbRWiMVw0sgbjEA2jFfOn335n7qp/gd77qx0vYjOWtT40OwwUmZmDx3Ch
gLHXgt2I/PlGAfFWLHK9QChf41ZhQLuXGtdAOuRny6PbAw6A54+bL5xQehM3NPLW
yvIZ4TvCGD100IG60WLgYcRAAI3e2YrioAATziBgZ+fkPEykOQVblTQ1Ds+3/aT2
9TPFHUDLt1kQ1egfSslPbVhx9fTmqCGdQgJapTovm/1cXZ+RRvl5td1OfhpH34dX
o9x9t35gyUlg5o4kdRqUjtD7GBdgIYIr/7NzSr+nkWodjGDQYiHUkFUOVUNzetvI
me5Sf8rRqFlivdcqvw0Y1TqPvVx7s7Zy6TRcKNFVA8PxopIrkHSey0KdpgDZpmIW
B1c8wa0ghqQ0pmWxTcCf5LJtRfSaXFc5o0nTtCyItsvaT0W1G2YHjTtMdyRNXAHH
+aWh+6/zeJ1oyhXx2xv+bX5nduaGyxcv6obtqMa/2RWymvUM1Qr9zYKvkaPkoLSg
bQOCARMijfU3fM/7YLC6hK2E925dH/9CY6GLFzV/N4YqELhQE4116uxPKhqSEOp7
hMhG02nicDf/P/aWYhIB1xiVcj/dh8AS/tZvAwi+afk+nFeiqAjh+ms/L72xSu/k
iUVvltxx40N4ODQ8N6+XC9i4eBx+x5SnBjKzTlOQP84fCf4OtINTVEs9+iT3oYqn
zxz10MKN4iommrqalW3g/jx5L3GCDE9z5I8wzn7ZtAe4KNGKQTiEOReO5XUty8+H
SkUuE981gbtcFNHI/tuPbkEIczXLIKgI74O9P+1XLn241KTQ1zeA31EhHUmyggUP
JC5y08uMyTFXdyayLOhyi+ZTHaa2GrhLxA931n1sGstoT36q80HTYRbOSSSJmJy5
PvQenXdKHiPSk3XNzcAzfzcp+KZiCG3ngV+BO6PqPUMfIlf/L8xknBqm3JcMx9pQ
jalB1LeNVR0xCyLEIKmeTcgjuxKLTWae9K+YzyhV+79wsG492PL/jL8SSoAa+bkG
CSPDiYUKE9MQaJEv5BzRCozXiuncil7W2GtgyhyYFKVnL4j7x1LJMhJgV9cgy0GW
GgcCcrftXqgcB7OPEWrqWxKbcj3EC0R9RlpCxDPH3RrKenCOOYjiQXzumVCrY9dY
raNmDCPtnXzvw0TjcTv+BgDfHXf/45WCsW08aod/Eo/gvBwVR+Qu27ruRV1rsGD/
bopghyk7JpW1T8G1yP1L4EZO2E1FxXYjQc8MzMaO/t4vJ5hxZF6UeuaaBM/WulOM
YlkuOHWZz/+GUjM4Hmpbt5JsIBmu+X+Mbwj8fuYUMZHZe3ZttlXuD7pzD1grGqgy
abN0Bm0x1bVobwuSeiJqkETulGFP4pOSnkADxouLARNikdQpvij+9XPZkjj+rgx7
K5EGjwoqhogULAYA7+JDRhDTiop6VZhdM/u/C5G4tsnM3YlCPJMlektFMq7GBg1P
gAx2it2VHM8ImSNY6bcVZGhkVdz3X/pvEDhTeNbgXYeQRmUxeNOB8mk4eVBcWq40
3RQ852ANa3oHXW2XsgOXvor1quQMYAhpTZ9LLjU6+u6nFYyrA8dUS7lDlKkJWTgC
8N21a+HcClaHWLxVKot/dshc6JiPAGxQroC9KBjrnOjGznaVBMDCyyR2zuaj+BmU
mcuSlIjC34deSLbeQHdKnPzswu9ApOGTnQ/AiNnpNf/dDd8GniY56Ph5MTPBLKRq
jluiIV/kFaLzPGM/yzs4S8y5SivJgaQ31HO1eCeVSYoMfGkveygbqkd9vmXcZFZC
E9919WEjGTg64kdh7aRBdVG20raMOw6l46yQF5aYIIG0vEUZmef/4kY1ZY5lqyZ2
OU2mnS2qMGu4rZ7UZoCWNf46v+8bMkuelu3Vj9vopNylN6GkM7s3h29mmF7HBgvl
e4Z9+vE2CKF+JTnmvWwlgCtR4oQ45HbJxLQXx2qhXOzY6Txk42FyD27ICPYEXcUc
hIuFNLoNiSYy4ukZAHhCDDuUfqY4tdUu0700NC3pnulSgJ2WzXq+AfolHxn9WnPy
y4VXaKy65esEVZw4hGUJHinxGPssA91QzC1If/YCoCfOWbjKO7GmBBu1OJTyB/cM
lT/3o39T8U/EZinZBj+OHESYzU51oyzcHprKnXhPn2dxHUx8xoF30rCDU9o49qco
iTT8dLpwuRIs+y1sMrmj1/dQF4vh2oEryFByvQrU8jMADapd9o81ZajP/MHQay/U
boYMnBPUUKnPa+dA0a5EkyK8blvnA1emWO1kbQXnLgKJHKO7eF50HuExNlOmVcu/
XyxFv5FAx8d6EzBGnEsQTl06eCCeKVQoJoE7iw1OMt2ft/rwatwtxQxW0XVd6TWT
SpjcK4qwIMyWCaP52tHsZL5KXpAfGBhNf5CQxcFM5SuXEu/GdAO4BUo73tIT9hbu
G6vFM3F912bvSbAWxQTc68vMaguqtGgjOi9JNF6/7D6CjOs9+398EdG4LT6eb0tZ
ZdAeIMIu0KG7I4sQr7usnKl23DJJpMbC4c8jxq+UJyd+Q4on46byKNDvum35c9rc
vU+VEkMH2b6PshZ02uBcbfu6aurNpU5p9FpE0/cF0COYeLAnPUwGsBx+4zPgt0MC
6zqeGJlU208cOFvV0uMW95jy0olDCv+0TW2ODT3yC3359/TphqDVFp6Ye/NXm1BP
KB71SvcHUjijv857Vj7WByjz0DBFKncIov1GLd9LbSo3wUAxQKO/Q3K4SKq/JbGq
sNYRgSoomMeCd4e+BD1HayaaJMhLhOrUr185Lr7BTjOO+ZN4Pj4jUJi+cKpEzB9W
2/JOWe5jUTBsNsl2975QQ5cvsS53q7OZRC7kB6kucAhTSV63PMc4ZPrDVteqKyeC
zRAy6c4Z3tVc3+XOggIzt+NlXm4ZOGcBoKF05pPOhl3anaWKeGmp6K237OhJ/CIm
k9gZeOi2FoogEgngKruF93my2PRT4etYjZ+pwRvrbCZhETprAJ4pcS9VOlp8iKnp
0NuXm/RrYABd4qx1ZEjPR0CxTmlXDcO64EjgA2nRp3u+yst1f0FXzYHfmsDCeH9p
1tXyVKMA00NSEkNoRJ8mNkG7ZVtF8X7ZbWyLLr2kkb+N6wjFgdIxrotmP3T9ooFD
NmT/LK1L5F95f04YzScOAgFAKs1n1rvwHWSzoC9QCiEL77+KEgYIip5unl6dO2qD
MBNKBaXalPcmLByzyoRBKPX2HghTH6yNeVPk8I7ijtSH4vI4L1Bn72DznnlTvq9W
BINfacrhFQMZVIRlF5wvZU15m/n2VZgFJk1R48vbrnNeWLyhXQtCDmYnF2zcyeyh
+QZTYGhDXm8N1r4dJqEYY245bVpfQVRjJK133Xz3QMgga0NyslHCX3ddVWk26r9R
8pTI+83XnkXtps0U81IQk8uMFDK6WgdqkJ0eEDyVhEulzrqkTmpaY9+7fvW/x8uU
aU8DogBwmFGOIUxrpS9I3Jpb+O/f/hWlFHwFaJl3LWqNknwBnGRyWzrmgRx832b2
Y6wGav3gEcIDyAgngv0kElPDkOhEM1WFl80dgZ3MMdXD0izuHh0ALbonh3jMZOag
+T2JMZO1NbZ+ZRRaxO2YDOHcC1ss96UHc65seOMbrIkrrnx5YAmYQ0ziIKr1pwdp
1dOA5NoMFhF+IMQo5JD+5lTpKadr41yWTrVWlsgcTkq5v6sjmrEAvvFG67mU96D2
cYjaabi0dcjstpnDZsIALCydUYltZxVqDKSN1BSheOzpOhwLYuXr/yIaXgxgGHcy
xGJjTuut0QFQ9jAJAN4s6n6K6lsfIzxLOC74G8qr0mn1fScNBy5s7SFOgzwqWhk8
rvR7Zh93aY8uY/Sg/VJhNq/s/R87nWCVuQT+/qBIfZfoyN7CA+/s8L/8x/EkETFr
lt3nnGTFcIwtLGJcdnBfGPeC6nKInSzbrQo1mvnbF7naO4SQxIyQg7CkgfNoxR/1
QhzuoDtX/N9vzynccxWY1UIdiR/zg11+eowVVkEET/7YByW1EFuhYAObgDBZcxsv
ZTBUiplqd+XvOoSZUUm+/BK+y+ijKAxpXMbH9wYiGI/0wffqKmxLVMRrcY7qGHp9
gq+agkuMmvTfBGlhdJkLiB1wi/rVcn5J4X5lxz8GA0a71A3EzumTjU/WKX8Zm2Tg
2EiD9NTh8dJF0ZXOzPCDrGGMKZbKEObsxBygK8sNdRVHkuRNFRWmP+RslUyU7MyZ
Vga6ycPN9Nf5JczR+ztM/BFHk9Y0Homfo3Zi1Wh7CN9+kjRKgPuBRbnfvOWLYGC4
f/G3G7dtdQWwdr1ZB52PydGFdEthntJkOpZbghdAeT/QHCR4UOCiRc3ZA+jt4dOm
9SqlmgDgax/42OZ4pyKmTo+ZRK541jDvnaJl4yMVfTTNxmfRWpbJ8OaUxsmANOGX
9croWIu2PBThhGRhRkQ048jomv8ihKI6NwYsjpQH4fFi0FUdMd7Cc+fXitfueN7N
IbzJPcATafYwDaYp1iFhDayxIddFBLL2W3VJr3YN1aKTiRFnaZhyife29Ywu/39Z
+m8RnofnCFTfJBX4S2o5+h2DNWSJsCUYRQ520J0iR2FHCDkq7UzYDty5Gu1nxmm5
lJpWMgCGTUJzPyxA/Zix7znz04CBqplC7XLTLu4VAlciEvKuuFLcLB9c9OvLZfFb
KZF9gWB4Lnk0xNKmqApsmIRhmgVZlX4pHkTrr7fwD4gMqwXEkg07yoFcOZisHVHM
KDOaeLzdU+4I2paMfSmvnZut4uKX51T4Zr/bYstk1M7shvre60AMJnsjxGeyzcx2
uSIizVJzrJGOvGKgpO74gA1b/QzwurCXsUvo0y9PuTPMYJx95xIA00otnR9A5FFo
p5xfOITYhV5OKDRgQ/1yDf+XJrRQPwXQGgS6LpQt4s9MhgX8ZCpK+zv6842SLLJx
LkaudrbN0/prYEAuTZ7mO/u273DE97sESqC60CP18LzJNws20556FAj36681PGTr
WMor/A8MpjTE+LsM1je3zCfi0o2iLSLnRQtwtOQB3gprkgr6/GQHxkTQA1h3ZNQL
unFHbotgU+t3lcYHyykBbT7ih0b35bSqvcq6HfCiUaL2Wq99r68LtLB5hL/Qz/su
GHWgAd11REFsR8Mt+LWaTZ7z8IqCWXynzVsa0UOGGxAzhbYRQFLHbAyrSMmFY7Ue
Pvsi3izz9uQ/rVDyKEEVB+snlROX/EcnXqGZYGG/jC7Kx3i60QjMAvLiQGh8wsYP
iQQiXP9WYxfTTgrJe+emTvY2n7497PKr4mmMAUZEOFXNKiARY9aShHT0vgL5804O
cBbVNzrM6pUkqDwPJsCnSpeIW9ah2PBOd0KN/ZC77yMKwT1LaEFKhWNFUNS7ocaQ
8y5J6c9+o6Hmqu6KXMAWZf12mDefxOCKiVG/ajQYu20hCbn7NhICy9XMw43K+ObZ
N1/SAMqLzXLNLmYRjz11dwtla17U8MAVwpiwXgs7T2SSA0TUYWGhm/oNKSdo8+jg
0T6sBK+IdQ9mxaqK7kXJ+GbC5m9dZakd3NFJmK+E3zRK5+bwyGOdVh3RlRqIFbYK
stOeX+hdeteXX/cDxK6JluGQkmwqHeIMEUWxoGxAusFoQZNR+M+PqqEFc6MtWxe+
XGyEYSjOu0t4qz3UmR6H3YXPxL3kkHdr1m7ro/CyRicRgqasrNzMNmDdwEvLbRHN
i/H5TCfX3k3p1O0TtAy+Jt0Be8OB5/TlmRcqL8X8iA7vEopdbrmPZNlEjZJuIRyb
3qCZeTHZkfje5wCsMO3a4S9eP19cwk0xjj0vKMHJycLezTxwZgWo+Qb81e6CNKnP
Xaecee6feB7oOZa+4/f60xGsC9kIfJDwxuk6nmKrtgMeecPHItlk58bMCr2gIhKA
VRkbsPpMQyDdRY8Mt6KBjGoLwj98kQpP/3jPM2AK3nLEIEDgHMpx4BTD+aiJz1OA
43Pv1YZTdIfb9yNKsF+QLiFBdb5ZcaIyE+avGkz42tsax7NDhSx367CW69TEc81m
+6zyKo1RKfP50LkQiEwl/iiJQW3xJ8xpB5t6ZMovUf+aImz7W5CM+W+QTXFNbNeO
haWbT9zTs7uEqbHBMliHKNeIx2H2AxdYBwMxASkJxT3ofzYbFJ35WAz86PMO96pL
lCqRAJfDd2kKHYWYW7v+ANbgHlAkflW6GqxGHGok6EDbftIY1EU2WHwTuIIpar8X
WjUzaYUAQtxrVzUjilp78qAy8eMHkGYsMDaQxDKrbqsP5Z1OJzIUpfjq0+iPEOdT
FBL4n47BXqn5LODfm2cVh9hNe8trlHQ/ryQo7dOIrPiAQqbFAdO7pVPqGdxWQZR2
SqLb4ggXY3a7/SwLkIdvbTUP8+yDZcFlc3gi6AlOBP9tkjjaVmuocEzIC/pyD+9c
H2oDPq5U0Kmg2lTubZnWIZ8brYFyZtygokDG7ZgFwvWzGj7sry6Fng9/JOdO3P+S
zMumyhkFhUlmYpuY5DHcFagJ/Hwcp/Knc7jFfpIxCp51sHI2B3jwExBgNtab/lQs
dPqBqdX+dJvOeamt/9lwKrIb59eUFq5Wa43bKHP3mXdh5GFcsTAY4AIzDcnwhyRD
2lkwv0MC0pug9fA3mK0OWhwIS+ZzifparCiEakckPjLgDOY4gcrHKsBLieBy4+ds
86oBU5ORjC6f/MUVsiVTR7ONsoLU0LIFa+EL8ky0wAFJCrKqL93XLkI/C/N6wSmp
S8IrLN0tKGO/GEIliAw7q66GBpmjyHvByI2Kx+m8NwtKbQJrjkVPVB16DL3OuAiV
0H+5ok5DdpRQIuAYdD4J59FqbbwfThqB7T66/lGWHzC6ejDf5JCJQk6Erauw1gFa
OdgnQqvaEwDTk8L/xTGmhSf36XOKnSPy6CFr9dT0EknfC1+zxdjKIwLb4+sWpIym
5avIMpHrb6y5SxnzxARbcFt/gFNzT7N14u9+5N4I82lh7lYeDmbEdzCWWOebsUAe
BQyeKw6gUk2dIVj/usDRQJ7gQkYqmKuBHcUaYTog91ylTcJarcKHc+7bySybBg4C
uH4bzJd8J2Xu/dHlQ7zAPiDagCNDLZMffTgnge0Dl7NT+d3sekVR11gfgLnqg9Kr
U9HDI4Yn02jtyK1HSEdbO1ZvpzmrZPizRC/qzcW3LlXR97cWTWGnpq5hCLpbpuEL
lHcoZNB0iEi1Jlg3z5jNpdRxfCqnuXMW8mg10ngUcAhonu/mycpW70MPfBVXk5U8
Bs4EUNE4J+vtdwWa0K0cyMQEM8jBlGv3F3V+N186Tal+T86OC8CGcuMPWYvNCy7k
/2+aY0C6jkXvXzmppcZQ7c6Keddt5sCyI1hPURS8m/9NGyK6kPPwJI8YcccIZHb8
ZMe68asafouD2k0GHTctZdXJfY5kiwrOALbYYzP1AErZi7Z6Is63aXnHS+egy0C0
gPvUagW/sa6vJTYZnB1PtXXCLRdvkkRkzKP4EVWk/VcJjG6pt/ae/omiUsfLDt1i
EDH2PlcMl2phs4d9simVeigHl/Fy+AB0x6VDMQwgWK70qqqLXIxIepu8jsqiHBCS
wn7T4wK+Johfq2K+KaOwjwoKFrS9KBO9o4vmPaW6adC+RWCC0OnfOs5DZef1Epri
U4X2lNUhfZ69ozXRtis7dI84Gn/MYfExwaoVCn+32FmtCJfVZK4nbXS9b6glZ9T1
lOB41tvAgQrJNU2UJ15hp/erFEFth7gZa3bORKWR5JqBsC5OrdC+klMVN1nStmGR
RUDEenssPumQITJPqx8ku6BA9+zO8p5+Cnlux31RaUr+8jfOnx0km0tq0Nd0yoKa
4g0ELqpAHCaAs6U7aERggN61Gdk7uWjLtAJg3hBgSA3I5Hf79dnyEBwQ+fmnvqK+
QIFliiiMrbnzBdbLKwW6enDw50gPaN2AC6xJeqGDW/0ykRYq4Mp6zpQqWflfegfd
m1itYImb4F7sXjEa2E9MHLUqzWbA2DorqfgH2XgfYAE1gs74J5RxxgzEvGnCy4X7
9RdR96oD0d2CCWM3iLBjK82Llg2Iw36eABPEwLvRCKoKs7WuTYHohC8u0hkhNnLL
ju8a+PBKMDnkv7ZWt7Ro8mizSdHSFyJBEYRJUqKr2GOglUeG/0LqbkJ1zhMzeB4i
WjfW2B/3HpHcaInKvRXyR83DHVchvKsm+HPY71CeHGxzPGzefT1HIc0YNXJo9Waw
Pt1Lib2Lz6KqSqf90+HIlnXcb/OriR6Lm41+vmAvakwigO+vv4sr8sqga2D6dP11
DbGNiX4bvtc4rJm7RZi5epRwmxnqHw7Dkn22XrRxzKdRo+yum1H2xF/XGxd7yP9S
svK+U/qJAi5r9xQtlPGG0EDxN61+DlwicEd/cE3yodj6NWNHWMlHfCTcXUWaql0N
M7N6ZQ0bj+V7iOkhaOetb5bW1fxG2tAkKZQYX5IcvymY32eWE5kouNQz2JQbJP0q
bR5W5O/stL1Ndh1yIQwLIHdi6Ofhm469/TkK80ushR3xqf/S0rAh2A8QAtZ+kBLM
AWjcD2CK1jetpiwiSib2OR7YT3KJeKIMfkVwGTVaZoskrmvs4fBI5cgEuoaTxvSx
oGkxHP2NERQ0Zg8LzBXbADINCKec/xw0zYTUAcs6F1DycKcUQnOeQEz6GkEMotha
cogI2oYdb0NZABoDPmPsFkBbayokfYjoif7l3tUWM2p5xaa9v8pTOwY12WcXzA6G
WzRkWUQslycjXyVCZFnH7kHrQcqHmr+s2892Wpch7SuyjJzm/0+hWRAoOsnpUyLG
WTyj8w6s/aFOD3cYJ2hkOpFnK2kJ2uw78V/IPwE76tfr5mGcAnsNstyCX5gTQWPo
w6+yRjIoTV8DWZtYYXwqvMKLJiAXwsMWqOVThW7kHIsBfUAKnH71fUqXr/Rljzbo
PloAzy7c2OTVffU31Wu3py/iLp1AVxIfoh+cX5OSWUgo0oL3rC2iMwxeESKqQdyf
SUV74/ggU/PHYzpFdJOsUCl/kVHv8BUiCNk8pWDXaWF49i5iUOCogoTgptQeZVV2
hhNsB7asMgJUXKDKK2TplMlOGz4RTmeelV+xJelgSDNvhijlVDeJsOimmhoqCiNW
r476dxUWIQo+BNk2LyoYyjpAODnk95YEk3RIbzn2MewdybSrnErU3IXTeWUuYWIw
+6gmdzbPMVIGHmidvVmGOWQoPypPSD7Ehifa4JzDOBOv91yl2SW/oDTqfY6DOYCJ
esvqnT/r4G+EsMu9QeVnp93+GLINVKDl7xCgB39uUpak5gj+58KcDiceS5+SxwuV
rxDfMh5/P8U32FJ5Nwej+bi7NugThlJdDjuL0fv/nac=
`pragma protect end_protected
