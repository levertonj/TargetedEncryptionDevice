// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1.1
// ALTERA_TIMESTAMP:Tue Jan 20 08:33:54 PST 2015
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NabY3FIuz4j+FLYevKpTyRX3EyhuMLq0fhPS4gAKN9DC7q3tRm6GhFsiUp69I2gA
VaqThzQifmLmXR+4WqRiw1GVnfypYrXhKIBB1tdWZF1IF7MCUMvGyCuwcP2wgMxF
n3WFH3mNeHStYbkxkE22yNcdj7vYw2k8QRkIwdw/CSg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12096)
8B86wu7vKAhb8K12ATKNaGDClrNeH6MJai8qmq4lZBNHfaerjF8oQnNTBzJrjSK4
FeHnEyi3n/mJ7CNSJDhQIAfs7pLUYsG+dCLQxVoyIWid6YR5qtiOWtLPDnuJ4jtO
rsL0GiTHGQCP0YJiUG6PTWUzR/McCUszX2OmJe5Uby3PjBOA+CPIgNWkdU2uqSVj
aC8qQ48sMzdcV2WRzOctlKy2DQmSaENu6tCw4aa4yKCuAeoBFmrXN0DH3/3q7C4F
qpk5WELnyL2mRF7Wu9AdjKhuayaZehhqYJuihd63mGJznOiUqjYIyS+1MzBxfEPr
RVAuNjJhnGT2KipqMMNhIkp/QSYhyHXnzzTYsPaORtYICAFp+jpIsP1jzfPnrA+5
Qht6l3esO3UL9h6L5e5j97McZXTTOJuSGmtK+pMEGev7tvD0q4dKJ3zpyqS9wsdP
bSyzhO3RY6SjWhm0OJrdvcaKBebe8MYd93LxGxH8FeYz/RSTbgIvg2z3dkRDsqMm
AkmsJjwPdjyvjBYiMY0k7WBSFPpFhN3EEdbfzRAg60o7P++h++tPrqoewhtDY/vB
FAy0m6eQl3wqSX62NdOEq6RIBQlvysNrIJsvgcLJtT1NoLR/UVf0/he/RlpuFPgg
9EkE0vQls9SqyRVlL8XAveqUm6h2bF8FQOflTgJLA/T0uYM34lvSse1WwCy1c8H0
Efq+Ud5KpTvNyIK5tvVUabBizlAJyI7nTQhvGrmVHfDtC4OjFu3Xy72ORRWkKj7/
m35j5r7xBS2YumbXBVUiNzGGKl/LUUfg1LgtR7c3LbK7wu5KuROF0StlOLFpkMIq
hEQK8dBUeBVp6ni2ziv+TvxH2rdPCBQ/7JlMBuzWTpDSwUyzTpDEH0rTOd3RAGqS
ighdIzJ2A4sJKPG03vNJlx9vmSR+LC31HlaUb1Pr1PSUT8q3yyIKuCqWhhgMBUbJ
s2azW8kWPRXcW71o43j5+jCJhByheN+T8eiOHU1z7QB+ra8ZEBc2+GsS9Xjf0rZc
p/I5pQeXFNXz1/Sl42HJniLAX2yjW3zSJh4rY2Sq+uXmmOrX2Mz1iLl1CnBJOi1P
LiRFJILvmfE7pLvhqyhuEkR9bUNMN+5cQx6nx1byc40ndPsiG+pBLBiUr46J/lSb
cvBIC890oD8J331R0lEmXkx/spHUcQhV1/zzd3R2lU13F0pveTnn3xA/DmLdLazY
kgWswiyFEjkQVwv0Y0rNHV5PMpe9ZYX1m5+qDqg8gHi95CH4kO3Juq6A7wWnemdy
v5nZ7fIgTsbhIrBg0WiCdCjPtCuouC47NJy6MrrJx3AJFZIdlayBlssMy1M58235
BM+qohSarD33FdyjJhmns/OBvkEvmPWRnvRI0Xs1Timo0fnbefbw0sCRNMa7LI3A
LvPu0w6Bf3UnexAEyc7Y7PK6xCFXUO9cBtWVQPVImkxK6mqYHkxV1cHlrBuQFtES
g5LIR52XEYMm6p3SPicwLjSzIRxIhvMfvyfPxnMVqiJUcbLWoWyvN/Hgp2rUBM3o
plkm7U3J+YGfZgX5XC14EqCgBovzIiWjk5mm4DzDfy4Dcpfhm+n+e5rgepxo76h7
UTJV5Lb5L+iyAegd3BVy+bRt6kXokSvBFKqUddz732ZmOfc3h7lX7dE/McGbV4K3
PWDX3JI2uQf3p+1db+e1V3X/JUNtrrk8IhwoUmnEZoftlDMv1vRsFmc7NOqYJBWv
OOzBjwJDeCP9UAEa/S3pMYzUKxpAhP9NJ14hd1agSxXK/8lLzaneKiAioBrGAi/E
Mw5uVAQLgwb2r12nA0Eh/BUekOy+Y46jCP5BheBq4gKYvjIq7oUjLcjoMZETBGb6
0b9JAGYNFQwCD7CrjcMwBCxYA/Ia5DJloz6FOGLd2C94OBgIdH1GOewCLn4JIJXq
GlgxMsRjGg7ZmjoX7Ja33a/MH19C7WrUVZ8GbHYP07LPesVEddWqaiMKWnhgwuLB
S0rNEQJ+AkLgsmvcKYWS+9inZyS2VNQI7TfGYVwCf6eIbAZbtmTK6DWCRlQeVGe5
esKvjcKi/DqFD+V60GvQ5PUUZfPdv6f7JoW6Pb9YVRb0UbB61yh0x/kjuXdo7e37
AMBEJqig+a8e+YNMgLkWCPx96XH3zz7XzXeZrr43gE2+sAcPbhCasoXSQh0PZj0K
G6fB0Ub785OMIbeWgKWYyer/nn7/fG5g7Gx6eH14D6Fu7R7v8vzxernO7pIWO0Jj
aqan5O0wMcbko6SX9j3kbQMzNndx4kNI8XI+P6K67AjvVY1Pu3Clv69Q/QIj+B3D
MlK7PMKFdokzJG9csbfyu61Sw/kKRkG4mKpZvRbdg2BLF/JDAwetHx8YQWRI8sE0
93vAtAzHcwx1/iAmSEEao9MKTSKVdclWVe7h/bFBsmJRv/wSRAV+sIk8zRY3Ds1s
wWvluk6brfI19mEMz7J8Xp+2UV+z6RFG4xZrWhTKluLmzFFtTlIE9FchKIoEJLKP
sGEPBYFn433ClUGMCESzUqXCaYLQSGxqbiPSC8oSSSqpqk+RO3Kk0WoR0NeZwl0P
9OcLSUcRth9qNmOLoWGhzloL47tn9z8mtocUDhYKImuo3uXTZQmLcQD8qSK+f523
NxcMVD7hgd9dH0Zs6NcwMIe4fiVdnaL5DIVvuVG/CFxa288mdz/xX9R050SwhB6A
hyIHg2ZBaHQ29zJ7EfahbbJXoMZDIvvhBk1VgbxleXnvOgo6KI7azNv09NqldKlA
9kQzz/H46kEBgZsIPUw5XOUsUYbflk4Bjd4GSwVEzjHF3wGp+2+LE2EwV3aHx5gb
VCOulMAPSogn4vzz/QrSuxoLUQjd1g/KnyQhsvE+Hsadv1mWR36OSllNy7hY606O
qsA0LmJiCnc19Og8GtIy1A4QLPceQXj7DjzhzFzzNls+2V2N9gdCNOYVtK62DWyf
53yuodRTfqYXEP1OmfsyifgoRcc+LTo+yJyUMaympR4m1d5AItFo1Rts/B991LBo
yIl1Ko0FrkdAUET3WKWTnwePc5uScPyd2vzfWdb0BuhXLmO8KXB87tMd/UGoqF60
PEPNUf7QFxPughW484bgoDUzlvcO9RB6ybRbTJKbZMMJgMqRsYKkgHctONaUdAk9
kKMQa9FYlgu611LXukMYEY+5xwDoWIXxLzLuYvB39+N/nQtEDSAaHh7+RJtSSdoK
fiwvP/s/12JrCpFfN7b2fWc7Pwe7zVaFnsVRwVvpB6PZByaVTe8mmL033EEbPMVL
3ri3AjIrFjuVRMFYmUxkvdMOxdWtlrB5vx3yIVYw66NoBDRorj1NUxDPb0UaUzvA
JUkxbDIu77KpFWC0kY9hET2CtUXp39GvQM+kr+BSSCgIWjvpg08Gu9tk6hv9XiYX
cuHIi96KI0kbexPyIQAWnu50hyegtdZ/WVNR8rFywilaDXKFhDfWngG26WSSdBli
MgLR/T7s8Z81humBxhcb3WoAhejVTXvVv1OkwCuzgmCh87s92qDx4R+3h2RQveJw
qO7O9hj3+c5bfAvfR77eM4mwpzqG2DRz7+hCaPHMgqNTIJMjJj3VhdRXDSp4OFOz
c0c04MAkHJ7gSVrzKxINEWozA/P8B6lLvGIxIj2+USJz1q9fvfXXFVvmhQC2su54
lRKYXyA68roNB9Jjq6znP49+C5K2WfQ/M083QHflsHHn/aHbJf58XmEi2TbBNnA2
2swQxKvpwkNIBEaSrvoiSPz+ebHKpbUaQcTxe7k2vu39fOkrgTXRbDAjdfe63bwG
3Z2uJwLkg9N2QPHS+lqLopetGcetCtIRMhfgYwFy0tIAreT7S7YQZXVlakgd4SyQ
XKuRNSTFpBCLeWnafXuGuTWBysNuuUwrzx8DDnM+spMBKTA6tvORAMUF0bz3XwF/
PD9Ps9oqX31Jf8MrFE7wogbywvINHeYGGcne9KsEY8/4Pt5yRvN9noPEqUbf+q8l
zEgh/saZSw+oYNhvnk/LRyZEycW30Pl0JlrbmLB6BFx0b8jiiwD94m1n382gtXIi
6Q+JeL9YYcWOv8edEtP8LYQusqn9nDPoZ4yIu2U2+7lxB9Hnxfh20yvFUz4HjpFa
5CD9j8eWn4EeDicN0omRe0fyy003/jMUetqKkpbYBK5pN/WpjAt5AsbxuHgS8wPg
pg2GiZsfXz6zbq8T8AyeuPiinSfqFzgXPb7NgaekwqnGHekL8/hUhjZ2xNQlbcxK
Mbs89LhmI3DYEdiVAnlxMYH02Ia3sD/laxTO5z998UjdQ6twky8T3VDvsTYWg3zD
w9300upjl+LfyERsF7d3Hb8/txBIGBSaYhzSj3la43OhSRja45PVfeK+XLs8uINn
XuxU7FnjrnNui3Jf0g2Bm/KdkGFDPFecicQwffmjL/hrsXE+bAHZiLDWe8ZNWdvi
Tk7psrbHdJPsC9UxksX6WuBYsPA/DIAk3JVnKHHerSapbcCTNLjYvOca9cRtKWea
gqS6e5RhsdrnxldqE0O0qN7sbVeczfsiFm/t1mcH+pMjzRShfox9MZeSyn4WvVDK
7Pz+46YVTMGel+FfOkzhlSvbce1OcobCpe1goCJMQQzDvr2RVEvcOYH15hkV8TjD
3pbLpzYr8vvT7kwyISW8XeA2QJ47dixNXIta+KGRkIcrHiZlATSolf972JoT48+r
ErhqjPkbrbPsyimpupcsZX1tzVaJfJAs5gaWHNNB5995IT6Ry+QpOsTj2ooQcXT9
F0E5C7OZrStEG9i6QSqaB7RST/LPEj3cMXlOxuE6hz6EKm12hbZ/thdfgKxxF0Ns
r6n+bOZw070Hef2ILYepnBE/RMIyirrFNgZTXhDgEvOSOHKbYFSvta79Bgkbbk+a
1YVGJyCQBnaRozwJTtFaZUX9OoY2e+oylx5zh7DGo3nSITfg6zOOMW6rucQ0w8YS
vsTLhCWnz4k/JxBAmWEb3P68/dzzx6qF2HFze6FyV56qJz9hb/LWVfjT3EtOglSw
xRZzPuFihaYDhDXCvupwcezME8Ulf8fO2z/Hfh2CyXsLaW59f/jsv5YqOLA0TGKB
FYgtY57ZPUmr7+zroU1jxB6Sbya2uLYyu8QE47KEazR//PCQPdNGra3J8RYI6KfY
6HLMhSNvw+BBjz2GJ5y0Wsiulu7HlDdYwzhWEj38UlLMZhS/PGa9fu1Lb/JGk3xr
OWGDCpjZfC5P3M7MpH9rGqCZaBxiwsIbtDPHQd3a7JQrIUgsGNymkCAZnf5E2foJ
GHxXKc8PeG0VsYYulin+EdRgUfcqTjuni1Txw7AZX9p+TbE4cNRj3Q+sB5aTAewq
XmKJmVHCa581q/JiWjGkItgp7ubVp3UH8rZgG9M5wX8/yLygWbekMpCOSbhYBCBn
OlInPHmmMd0F4wa6k1uFUHS73MW1eLfi9botYrhmM3bdlA2tLIlLzHwVRTfxxr3D
gz+6iRApkGSqVvnLtQMQZE4X2VhrHHE7BP37dWK6bfvPI4J0d+pfAjTtDNZQm4ht
V8w1MPp/2UcbF2D85BeEZVEpNLKzC3iezAL5hvfS1ySxmY426TpSy2iPJ1VXs3pD
fTYZAAGM+XBlRVnn/jans57KrS38ckD53/LY9KWlm1YPOUm0OnWmvOXBMz31yjBI
+a91vYAPdiMvJvkkMHuwFJFddUJMFzVCE0Mzra8hoXQosdTxkzTR6enY2kbSth70
edvpe796Ju2v4GHOP3iik5ug4v8jpwmeSMXv+yrmt2yilWfoWpuK31LFRQRSRSDZ
md/P4Z6q9hmHvwgzYsAFCEF12d5/G39dRvB8bsw07lkVS+C8wubdUoRH+eDVhFry
/icBYzFJGgfZKMYPaikXhCa1WzPeuZPkA6TMFCNoSm42WZMSb5pk+d7O+kK4tnR7
jJU+LgF3s1xt/fuhRFPUxO3Ex+QHLirPbEjdEqPAnZCK4EYJBqL3vg7MKtmmf4hy
k7d5XH4TWqVMT/VxEQYFKFujzO4myrzh4ZTocchssm6eNyFjbCBVhedcbIK/poM+
iYwQIOch4ZgZlcrWYa8golophxYG3yCzRC2k4gpQI94MP+LfhKYq9xYFP0xKb2Oz
OQAMmBTbfZO4dH3e+UjSiOQAbaKHopvnBOOinwunXQm4YnFVrGfv8o+1yqz+fR4T
XQR8uj3cSPldnyN9sbhiAjDKJFllOITcny6lFPmtIAJvGoYx1Po8Q8w2Cf5GAe37
qgHZ0BDGo9qPbBRTcX965Q1JWNb+lC9dr6Zq4u1F1WvKe4D8icBlFiEjlZfQncB5
2seBvuxnH50k9Xufz9OFD4DIWmYTm6+Z4EXipNYmSMnWd3lfT7U+e/vYQTlSgiyQ
wdiEFfhteF0xmedu+isE1MxfmdDTVLv2ZKX2m6kwtYLoiMtqxvNb4SFrD6rWLblr
/V9p17LQ0k088DN0sNcbmZ8A6yx9WE8jPmposp7tokdAPtEGm4q9llvisaCzoBAW
2gw5HfC50oiavVcAeWvOelMChyVhoEFVcR9Z5y6h3TvHRzgWRcaJgV0TPM8LMD/6
F96q3EfCqEJ6sTis3g9Ba7cjYzleCcY0HvKFk3lE+jnffQ4xwO7Si2S/o/IX1CeT
TzYkQalfJC+4+N9jbAJ0E/QONtPD2WcllytzRFq9r64KpEkkep5/J234lIbf4dU6
ReRmENPCeAc78z/hzSgJRdeilNZ4U3PGbM4CrnSRMmhYYGRhbMJ7dxqRwSc/3HHO
mvjiqiLPauFTBr3QWZogCYprbxpQHa+Namhs9K6oSb7QaBNcaAUa0R1T/gel7rCv
Vsu7KNXo2CNBeU/j7iiaApDfRszCxYqut/h3MhkUt78rBdKQReXFxMx2f1rdQ+RO
wb9WfzX0r0eBuaEEzzuvTxvutuODFv57ofj7WdOk8voynB2LcmB2BXDtGmY8vLOJ
Msuc1VzZlp4dO3QT7EHU/6d3NcLStX73oivbLxidw9+77FCL5OUGh0qddM7Xie5K
ureWrORpJmfAlUa//viVzlIIzki3BoOnVm4YA/lLwo7W5fn9BCAUKBVt/xmud4vp
evcChhHr4/OMwaHARZbWWfkVHXM1nsJ2clWe1dav12YFtTUxz9dL10Gi6buP6LgZ
FfhSFa712Ucvw5xORFcsU9Qw8KuLTJkHu8VySueWGNSW8FbIDagtnBVWGcvt2ib1
L1x9VGo9SrzeyURXE40CYRRJ+psA4zUw8DzGnZfmVGt/xIJ6pPJS1y33FBoTg1C5
eBCf2MVYynwIL+vzdR6lNkkXKB9TQzWAKUrHERxQuG/s8dsDb2ZmgFmMPXQv//w7
grZxDhEkdE7KxKOjTUMVg5L7YE9Zs+Zhlmcr+h5TSE4/cax8rWqpjzQPOnlCkoO6
NpM5awUuacqIvuGsGp5eAPBV66Hx05ovWiryTuK6zjHI6PGJodFnejE2zFo68hT9
An3BXqHKLWSbvLTLpxpGHYZcAwnmczaPTHjW8WVt1podi8r7lFk9e2drDeePgxMF
M5iTvfga/8iYMOIoQBf5Zxf5z1Ompjjh5CpupE3UIr6ANQocEsXKIL/XTWnZXd6N
qZlZgYzMG8LnUIJyqFuKEnF8OeiMLzSzETGs8mqOb9R0Tmt0M99xnpYq35h7FeDK
N0o8D3u1vxx+w/6iJKM1pKcqU2HolAeUKyVVUDNI1ioOSnqxYHKsbERUJCCgQcU5
Sfx1AhCA++Ti2qWoYituJl3vyGhxLQYx3iGtWcYaYPdF40yID90I32naaX5uxKPA
imCwnbbb8K023n6eip74Z/dxt4XYYCh7JVoNIgGa+tkSebjAssyvFtk4YRYvm2Bp
SNNspvgNP9P/mVMOIW+a7GvIDoNJE7d4rfYR8GgTplmz+AKYKADikbOnuu2UJi5D
Zu7Wn4+++j7Df9QmApQE9imVQNy38Q8sDUh7uQAyR6k/bj8OYyI53uGL3O6t69O7
HasZUHjYTXqAyQvCIdK5xw/5z0YYu0w64cUW6zFk3ytA7kPLTa0oVqPIX+N6AE9b
mWUa1zdLFMAbUjqn2tvXXgOQAQ7bq9vuE9KEb+ttBPm91nkIpGctYvVDiq8yUKQu
IzPtZ0C1p8n5fQGhilJxKz4zwj4pJh25zYMbizrOC4BsP5b2pPIJnySwokP5k6JS
rKdtsr9QyDlBEsLgSa8te4NK7w23fu0Eg4HE2NQwx8geSkCy42xCaYSOhBbVwh1n
DS3b6hd18G5h12kS1pM5Q91xGh06Lt8jWh5mJfHvy8DQGBqLEgEcH0b9bfd3zmhR
sSQ2rxZVkvnIqRLDO3itd6BgzHrWo84t2t8dYtDy/pkxe3D/gIQUhyxcg7P1htZ0
jNK19ZCrEOlrns2yHnctuEl6XOYvW15j86HsLbydDzHcLFo1bpXq59BMbHeImGoV
qe1wjW0UsgqdmfzlTgkqRc2tiT76hSeOIBLh2dSlBstVf8WUR1ikEWgGHFoGvHgA
/K0CnUe4ONZhs82aB4gCpU+dMXkQWvHOwp0ybLS1zw1eZ8vTvuQrZK4zi4eFz+X+
0F8JbMya2IsMMz3MElYLRpO6vo/2J00hkMH9p5SUFwC+92QbomexC8mDIiBA/enp
zVxDTKS5pslSQgb2zRRuhagmj8OavqofzdBQm4SzX+c38sgC+EA4xiaAPjfxdfpZ
Rfmy4yC2U2it3cRjlaJPzH+ECzoVNXloO0wX6SRX9Kvy9u2uYXrxjueEe7uEeubX
1TPyNOHQFSS2DB6xxkCm4wNYRxBPO39YErKCWdtsZtemQ7SHPEQB84FT6ygkaYfL
VCGoCIFtZx9r6/cGALlNZPu8iMQ5++mUD0Qi+nw0GlpK9FDdoXRE3M5Hyz+slnF9
9yItpjc+eh1bFPAKnYhlq0+SHrbj7gy8UIHh6z0EWYThfhp3buRbu4ImPoi01LY8
TQ4j0iNUTqN5UF7CglaJccKOOiNsTzGyVgOehoDGW0BEPVsXxv0BqBA+9l+seri8
3IY5f9JV7ltOJPRXUJmZeJa1TxJT+aTY0wapIKz6pz4l3c+EUeUoRG+PPtm7Q5dR
frUpoDQ16la5zDuPU0AEGQ2FScd/uElk/htMYNOhVDEN73m2fxU2UxX/SWr3mQAH
prCAOybbc2JGClEeDc93/y7gL64y2q2swCDxRzbSKtALmd93tHRkerKH2Imml8V4
v5Paxt7zX5pPzlqpX/zTziYUe3EmXbEgv3aAIwS9pGLDPuzF/9QLxn56mczswJka
hmG7k+h5jQEyzozzAbecdxv6qRjT0b2AWdf23O3HW44CojVJ4WaSvXcWHdQjKw4t
t2G6OSVPJ2u1hJaJhB3+BxJuWRKXfzgZZZjJZCczpP2i14BIwiX+GBEHzpEKVRbm
kOSIfD0TYOhxSqlPYfKE/WcSVSSRiF/qv75FKxBmAIBLx5C3kkz2lFblShk8cUFS
nE3I4Lg8LPhkNIJ9ACn9SSkhJ/EJ9NnJqNgzN6s9J1+HFoqUArbTRAxOlRLJcyUi
PiP8L8zVDtcv8Ba3A879kvjosN5Wd/4fnvbV/r0ulf2VfIKSwF8Bt1/873Yk/66g
cSLeWEngFArdDpyoLnPcIcKpE1GsqwudDjzCqYcxKIvyWFCFy77dN2wBOUpy3DU/
X63zzD0DDT1TMiYGBjRuIsBxZtZmCaHzFqeoP/p8L5ST/BFHPiOsq1+uEl6L+jgX
Iqc19yW6B13YPtbMPeG+xsWLvu0OvAgNclZfF8m2SzkrhwSrbjdid8XKKw12BJ7I
LEJxMA+uBAhdThR5ART4MAVS2S4mzt+2fb03nMrvSmsugVjJWYuFKkNexvQjYqr7
GArdfk+/1vUFaWG30qgGl5bi+XfPmosH/STu/aiu4rZBKzr4gSn11M99g8fgurpL
nqndJknaALvrGrdtk5yKmwfhH2EtgN4KKrMd6TZEMkUQoDluBqN2+3fa4VVgUjca
WZKsJcMrbKMhREYhetd0GK189yUWFBe8mSpjpD4/viofmntNTTAEXpshT2HCwpZK
hY8Kj4go8TVL0ieB0dA++1hK9jaVM4LrsBFH9H9D94xY+xz0yhQ3eC/V0doSz43V
Vgk3WwnYCzOXgqSFt0Pk6J2YUxsTkx26TIIlvBN5w3taHUZgipJ0C6iXarT7QlDE
HvIXch4dwjB26G6CjDqKMJWxsp/in9QbYTHOdq9cfS6HAkRO25rUBRfDnlb0qiWN
xbHp10l2zmbZwKYZYCBUJbGuMB2qP32M0qWWD6F6KI2gHD2Yn9CfBvM/1S3Hf+Py
2EHQXVxxRnsCdYwv/u8lv0jFG0jBqxRJZTKcp2qxm2UYHbj2pEsEaTBspC9P5jsp
QQAk3J0QsiaS9pgz+Oe19wi12EDig/b+H5m7SwV6cyHuidu9FbnZ5T8C5ODM3ZWx
p5pYEpSwisKlwz5QEl/+P3uOhOpYj56fcMOa6YKypwlKvTJ7s5Tt4vyo7YRNaq+j
mL1LIK2+9A4eeVabdQTAUZiyo31xUMs/UbkecnuiOm707gN+5q/wXjH664tSO2It
KZrZdo++AJN4Z5qogfRC+Ac8sKFfEeup8tCg/tLOfGdftwNcIPIr9Qz/xAkn/+Rm
GxN06nE2PMdglcC5yRcEO98ToZYcp0GN7sNygJvdy+/Cogsow8QtRapFNMIlQNe0
qHLbE8KIzvh0Vbtzlx9J9jow9iYTERYWgnG3yfdmvpkDiuCeKKfrSYvHN15vTvz2
FlG93LgJDm3zobDDjJu/JDTm28D1s9YGNXB6mF5GpxLIWtVMJ3tEJp8Pcezua1oQ
lW5t3+b2hX8jfDR2OoitXNNcdZknwIodZ64DI58Gn8xDaEG9+6pkfumEEZx+p0oE
JVQ/LOfhTfhJN65QqPNVmd/Tfjs55zScL4pBhh/XO29XUKQ5XLRMtxmd49km/cFm
TBkYiuQFiw+HedGAsEoB6JQK6395RfzJmZEFY44apDu+/jpJihifWyv17xwOfc8O
mx+pn3rTi71/bDIWKdCV5iB+BJ30AiaUHQklnFgbQ0VQ6Gui5TIDtxasB+w/XJuu
0LXvueJktr3p1LvhHN33ZBk3iTCu8s5U7PnV4wEhHBkNvy36ClwbM/r6CiRj7TIB
Qi5GnGPUar42ka2/gjouMEQwiwzoBjcuv9ooT3z3EH9Z0IzuaB3PUZBjxQEWfvD/
PlGRoXGVhlNi2vh6k+X5IU2H1OtnuJ4Q2LGqcHz16l9i+876vIpNHaBv5jjCobOL
+axLZTNp6QmmI6S/tDqgA3HMXohtEMdfGqdjmG8zyXt6DDHfOOd/0X3wZqxAGYVp
jWMgRkoeCDaHgWVHfe55fBJ7CzYHMTwJqp0xUsztzaVVXK+Q537Zj40SEPu+andk
OsycqpUlCOSBK8/ijT3K4uvl2WQb80k4mlWgfHVRuxUMhAy2eOk5Ae6d2rp6cNLr
gvnfLbxzKSpLqkz/FkmXVZkz0FdOT5V6tYq5rhcLtDMH/E5Of0yCRbB8VBdM0df6
r9l0HQ1Qm4jOVIAoC5S8fJWR6IEVydpYGEt01GLgQz9t9BokHNstNxPR2wY+kl7m
RGW1MVjsNWRIZ7drRzKuR8NvtUG2BiA2DOeQmWlm1YFwl9rfQDGmfFpu3DyndzT6
zoawhiqdWRl9MZC5wHFaJPL1v/CHm93ms5/KOrZ5ibJHgquURnOMkQ1WzIGbebcl
JQEDOj+NiH8X97eKNrR6PUGOtSlab7ffElIzMDq5FDs61e3nhFDnSf1RVffTIkvF
ysn4E2XvjDzm+x6hzPAk8N9Sc7uvFGY2Wlq1G3T6+AP/FzOJVYlS2bNSDabjNwbS
tDrVeZqZyTpk9g5pWhvqd6MhQze+xYhcqE8Sa4aQzs2hE7FkP+2mzAAyTQkoZfWQ
9bibhvlOQkfLe16ZC1C6VA2pIYnsknSfulzJVb+bUABCNwcQJRCVcxSs/EAMwO7D
AAVv6LWqOksOpYNe2G31ajdKb86QtTfPfonCTDsRnW3WBKIEMKaqFzZ0qs2KPPgr
NQn5ZXQEexqc0q3UUWX0ZneOUIoghxJg73b26xXJ6bCSMkcBzKi/Ft1hiQZt/zrb
leTP3BdzpIx5WdvCpo4qSoa1+OuvUSyt/hO0AarWYAwoehxA7dAriUdG3aRyYcfD
/ZDGCXMB69zH3NAXz+JXsPudM1kg30TUcZuD2kgknvN/x+13/4IG2G87wK52cLO2
pM606vzNhpi24y/GVizIxSNgdZ35MGgH+/ZFuhD4MVibnVuGJ2j+WC62WtaLNJvL
kjMwXmP9bmwyeBRZG9pb4btUIAX7PumVrKOSkSOt4T3vHZlEZEvgHwyXRijl9WiC
Hx+DCzpJK5LmL8WJ094jfM8S143vODRk+nPbuTDoUPRZ95tGYCevOQngvIYme3sz
fBHIFEKu5z4u2Rt5nXDRJSp58LI0XCmNl3iyvsJOLuuh8fEsyBMEJuaEolUpU3sQ
VBSGC76blJFtrKuGtkBx+xXtFmG8bAhoE22MMhV2dHTQ0rCj3r+9Hz1WuS7gIkUU
yfohWSUfTbmtq/tIlTgPT1fPZ79RdS0c0dRVZxC5MafZTdHYWpTGzsBWE5jWKvwz
0+RaUDMpDiwn9Up+9K2ZjXesIxn2mjT+v6sUUFW50SOfe3cW0HR+IaDtGxvkevUz
aunEgSoEzdLXVNCGsAZ2/aEtQMcWNS0O/8oUpkkF1k0KgyiEhIQlxHWVsEAD2LnY
VEQeqxlBFXG4pDKZIh7+OTgNeFTLWA5g3aD4J61nrbeyyQsWvm7i7LtoUFsmLBVS
0YeIauskRoZgxeZU7mtePUjEOdOklD2KA9iSvBRHBtsMTo4T97M/QWajOMqIpl9G
LtO0+dbSL5QKHD4NH4iD0SnJemMV6SFJZhAd/HHqfxK6jXxVCsiG2UO2AXPtVcVi
ZfQ8ra3vXNcCdaX0U8rV1oqDHeEyivv52yeeE8Qrd2XJ2mezadk2qvk74CBeGoEu
Vrp3Dus9dliw1Ugv6Is0lDqjnWj8GoMcTXZrUyp6bGoQYH4Ixr6ZcG1jImaAr9yZ
CO3wamrGzYIAUD0bU5HvNF4q7rkhQG35ZXIh3vlmb02d1wLHyrj/ZdioRBWYTCXW
RM2Nm8lN3Nit3qaKY3X7rjZbiSBFiBWX+Yd31HAsP4Qo4e/g54VG9tO3pRdo8lAV
GUoNAD30dNNvh/iOZpaXPo2eSANVKvQp7WlpK6f/i20wVqeIS1Y0QP9R5vdSsppf
7C0euyT7LLFJJ/V6PBtby8IrcLKbWT9FkKj2yzZR7zGFrlPFu3q1S1xD4524TSI0
aPBhZ/8w2oQxrjqMCPlt3JZwxboVO/YXt9ia3Qs+J//M1AVt21hCcfX6B72TZv1F
ffq/x45X1lae1pFbfX4/GQ7lNuKiXfXpc+3oUOUHXoSBLMXROg0LsoqgrpWFX7Qr
iGqSOb/zKQXoTzCdM5KODO3KohCxoeiSiNUZ++pYhwT9IUHGRlwT/ao6eDa9k7DX
DQmzwb6ZZyIbqAPK6xrVjC1W8nLsisqO4CPK7ZlETVtJTOhdECN5pCQzqFJFmgeD
/UMo3cXhwnfBzjzsBCOCuwztWiLRthd71c6rchGHiVfSvg3dc9aK0yDEomj481hI
sqjzAuhKA4JAXj18C/mxLhfyMGCzVydllvO2Hh+XMGfESN2/F9fXnv55aK5FvpY7
cQtPsqlEC23dGu/wQOjHtKdGsnhjOWB+0kWq4HewybOsi5AbrtM81OCns8L04eZa
Ht+rQJzdNeX8r829xnDRadGGXyhE9fg54qTcN/4ohAJdqAwuVl92HTGsEVq9MekB
6jzRxpLMSjONVjQgIO6VO3Yg4p8w9tz1X/FTWdFvWgonGAxdgQJa53jCi3YbeS1h
KTurxko+IBiW3RYpow9guCGRF0fo/u2/tAfwREbk/pJzNOP6uDkQ2/BP/2W/+5iQ
zJwyFuFrNnFwVv/4BnjOpD8MzJtxe7vE4/LmV9lpqCK1rGhsP7EEV6cJrO4iNRqh
ilk6clyWpkwcpHdhm9YlrwMY1vAaY14ID++srQVjf/VWub0EPWS/E20Tyhw04AgJ
EeTMFB/tJoFefy6ftNyB6XkbfIwwM+fxwrNDZnbVU+FusN+qaqAA7nesbUqeq6aS
qb8IliohgJwBRkDCwxO9gx1q5XBjckwjtXroexP6y8cqwkg43DwWIttLo1k5tfA+
XZWowFFCMFdmMPciUZTohA0RxAcqeLQJlM6ToDmYtqBt3Krkl7xttERUba4CMFGe
d3cbYwsgLl/mPSKIFQo0hzW7qINfXkTbxt3r2+2KZ8qPBrSSHB2rawTvIkXSnQyk
haxRDdptilEDnK3/q920W/8fQ29uop2YEblF1mxafxuV7nk0HDVfGoUoyvWL1v6q
In+zA8docFbcezKBqrCGg8rEt6skECzWME06FLrLZ0KWK8ENaHC612q1HS2vOWbp
2QNeq47e6R8rY4R4YzgoKjDZ5TlVm2/m1To+zHwe5qh+lokahtrd+rcMCyn6YiUe
FNYYbv5k2kFy87PCEMZzp+voyJHPky2FTeaFkztuhT1nrkLJECrBoCJ95LL99hBF
yjxs+Zy+fFY6dmOx5DDvCYVq0E690JpkmT/ZZ9u272rV0dyL61BteEOEgTQHWDEU
XJbHsKlxFg3Xu20TNnMorZd6RWoeW/iqUIfE3qtqXKL/nMuId9aVPjx48tIDweXd
oitzzK85gK5IIUCXAPz08Fyfe8EkyqwNyLEtZrRme3xZD1wTFLqcoiVdoAxw6lJd
OFnnosgQhLIwCY3Yc426N3uLEXRyExbUplxxdc7DvdxNWp1ae2NJnpk/q1v1++G+
uleJOD/u3yaKCavq1bh5YHYzhFVTnbrYbw2zD5P1F3NTUfrovZcsRBMtfAV1Lv+m
R8Ak4t4ZrjtTFIjo6rvkBEATImMsGoTj3hlf6ZJ/lsFyXK0pmLtOFs3UvxRFe/GG
L01sjpoP4Q6m0vRqhG1QN7fupv5VYNVXCbf7eS8Lz9Oe0KgBuhGCjSdFCNk3eW3B
SLpoVYTBaFeFqn0cG9OyMOc4MxDmPaprwUxTmcALb0jgZH6drvyufo2FXEhY/cGu
r9+P6v+lP477/r/XLzxo7/WInuDIEhTli9EgEFvnpbl9hC8g6PeoI7Qz9gYY/EIE
1qZzykVY1dZQzIsan4LbVMlVL9MpxEmr+gUjbCL9I33uEiaoGyuhRd5PlyyPgemP
rd5x5y1hKUvStqMEf12G829/tVUMg5jjQ8iKf1D2BQcaICI8Z6TS1FVaq4C4i9ik
Tu3XiGtW25a8Za0kWS9ixApOTYREVwyFpCtmUEKSHd/skD/+SwBoFfc72OXAqsRK
/m9vNz/CIOl2VeRkXbHup9wRe9HANs8reopQ6tL3HPgt/HS7IuY00FgnhtwJEJYM
pGDtnVV5Zuy3E696f/6eH9k8cYAYO1/JXz5pfGfYJKng6dwR3vTcuMfIAnJCPE9A
1a+1f76ypHyoUdwlykhLImNMDEC/HW92ElDZDIo7FFNyOwrGH2HjyqxscFAdH41y
LdwBgQw4s1VfaD66C2TB+pix4FJmRfcK+xsH8uHiOUv5J1iVTpgicXFOehTwWZMZ
/2fvgVcvsaxCkBRFEceZpzD7bFOmjOmHEJdvvomBmuAYAP2wZRzgzuTqouQQV8Y9
D4McSjgiN+ZpfTAUaOd43kMm8bjVMLdBXWtcSq8bMZxXcDiCnxSIOUAj37xzojyb
S8n84CHwccUDiaRi8bLVNEhKNTRc3s+/nke2GWoeImageeHlTkE3VLph/MH8dOVA
MbdPcFI93vDsK5rF5n8jerkyamRwpnp8QKo4IENTzM9zUYCKX0S0bSc/Q0Ey/sbz
ikL0gN8RQECfZ3XCLxW5hhipXJ0Zl6i6vPMW1YJbfkgKbo3lA6K79qwGOA0HlvWX
FkaChPUm6kilRUTwQsWH7TlOVbvaz85h7cn7Lh7GqjKlhsfTDiZ2yt88BdPDus+F
FCxtY/ygJEVHm+sGV0mgoUOiN++GtPL7dIEaNVviSuKVprl/fCG7yvJOBJW6xOUQ
vMqvU1haNLSWlsyUHenMwFpnmxQpRkfUME1zdj9JdKWkdCam2wmKIycb0VEzUmu/
ItWytmCVX7/0Y1DAk8QLKRXSBTEIdu6SIE1M8SSoOKBd7FtTfw6P49IirpdRzh3b
`pragma protect end_protected
