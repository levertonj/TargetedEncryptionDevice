// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1.1
// ALTERA_TIMESTAMP:Tue Jan 20 08:33:54 PST 2015
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cjLmb+Vk+JVibXhdkz/bAHU2paS2bjDfdhUnRisrWLl4EOshpohbpV2CM4fQYa3h
4E50GxC1F3+xV4ge3xENTw7YH/WzVXMLaxPASX9QpmenhS4HHwIyCAJHfdAo6dZn
54hgQFe4j/QeDnUVJ2vr5e/rQglIFuhCleR2AXsZm9g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13968)
L6kh6TsXpfKerI3L2jnSsGo0E9WipBIKZpWP2pUl6wQPfP8+GpAHRpe9S/DBGd4t
6mmo6zWov75ho1UMRwEamW4v1a7ivg56eheVQcdt8yiBW1fNUrOcSvl+IhDcVo0O
H6jhW0asmWnkYWo2azdQaxh9V/5Y/gALnGoG2UPpAdsMPxvc0QjvtDVL6fIbdwcB
6DoRPWgIg9ekO9daGprptwmao1cpAtbOa6EY5e9/jtgZSvCcD2H07+vgfYixlX4l
LFfLH2IIo0KIXOPvNtemFEYk6xYRRmbXYwu1wiYBSijXtk8xlAG9TK5P+2M+7Eiq
NQsnxRMQZSCtojom20kIaEs910D7qs1Vi1p6v38Bm0Llcv9M3MW4iK35cEWz2s3F
Ue/s/G+Gvr7ulejQp+7SkMijlYxiQ+toCZIL9hLpSJwBGuawisHQdaXYgIda8cfg
b9eUfxTIUlOX4As8H5Ji4mMQC1p9OrAPA2Kh5RsB8TiZGzXmphqnHBMjH4WfA5t4
jWX3l92AQa1TY8is2NQxle8TjnWPBkLevNiEiu1WS8RvRs+IXPajS3+7xrr3r995
kfj/HcM4lEtwiIwaKxYkj8bv82FggrUY9B5+OObQp6WXPXRBaZZVTf1aCcDPAZsY
Ku6rNSXyLRjukF1TVJzUhlW6ZGfhwTuC7wLk9C6aG3nNErRcsKCbdmtdKsz5MqF3
+6mCoU7+rBxWNtkQqO/+zisEycAn8r/WUSl949Cg82nAUJr9IZjkEL9VHrqvUcQT
yqORjSQa+nX4gAtIG9/rcuhpTSSoW3iyzbEAbtI602fwZu+1Jqqal0K7ZLzPhMkM
9WKduCQ/wOBuRqlQ+jguZtLDWUXEJg1eNW+kGta2UqoQzvMr5nP6QOND/zLn1LWF
NlzPZbEESmKALnwF3kzEin3wdNtprqrnwWkbuML5a4VtETI9FmjQp1PrZV3zqY6s
PTCBLgpitpEEzgLNFYmAc5hqt1V99PmslGl++WhITUWYfS1p+4tknz4Fz2RYockf
fOLpKUo2iIiMZGm2Pn1rhpj30myVYGlRxk3uLWKT47FlsWoPdy9kwZ8zQU0bWxq+
Oijr/ZBlrBu5tKH0LqYRgzbCiX+Gbzy1IRKsV+eYGZslOpclf6befGZHrdvbOEqO
XUoGGEr/a4by+NtnQWABvG80eSiegt5dpGeKWMZrlSUS/RR9IZk6gAhZgnmT/zM5
eJeXbBplYwCA5/Z6KKenIFD4m7g5jqAnZcXpIS57n7a1ramBYpUynlBkht+zvcTJ
ge4CfPQx+1Gm8J5I9PJOPLrKEnZakNbF7Nx1nx6Cbmv73Xt3jsZkJhVNjifwV7OW
qDIHvfJDNKzrXCqPs7ALbOERHyD3V4pf0zr+5UnccIn3vJ8q+kkJ0/Iduv3bFp7W
wHm0OyXJeIEgbiOl2YIDOv4YOhw52OpT7CjD/6dmDjX3qddX2qKqMuyica2G5nlZ
pAOjgpjWZaRq4+goAs1dsBw7QNpsecMG6wc82IO8x+kzKqeZu8W3RPRYyw0a0cCM
JR8wjEP2PwcIXCwjI/7TP245W+5jjazx9yeAE/crpxUB2d/B4HdFgwrgE5Bl/fUB
h+2RPSr48F6G5xqt4BwKDb5seK2bk/kn4MHo7thWPZUcubiNxtXPkCja4d2Mu/P2
t1NyCooSxQQ6eoeAzilisE3JpM2Rxy6LozN8hY75UfJ1lv3x2+iksXHw+qXtShgM
Zn+d51CVB7hkBU+94RvvSbl6ky5xxkiAEQ7WCH6VZCuzPoz3oui36zIMYOdLaHC4
YA/oU0qMqottPrbyYwuhVLqC5Jhu2/EVIGaAVYNIfzQPikLwDfOt7xo3566s3hCI
FT1jk3Anin7FDf7dbSzwA51/rzXWmQpjbB+UcELJBdo121CaYJTp74UWe5Y6SaCm
4zpXwQCrK9voHzKWNZdrPzVpWiZMSBJOL/4/FvlTaigDaHZRywi1NHguL+mZ9+nL
WtDWb3SsQFLmq2tVf665JPXkm6QoXFrUm3cL1P+ysAWRUUcL2lhy7JFHXA5SlsMZ
oeC67fJ0E8omyvd5AO+i6Vd+AyAxOEtCLjtwTejRb7WY1iR93ymPEE6TMZ7/ywbF
eU1QXpaPwkiwRbNU9MqU5HiJ+qW1iaZUgfTSyXCKdzFJwESpozEZlyKJ6hyxtDE3
LD0858WYTJZa0b3I4VEp70XJkmUqjf1KXGVmr2rV1mWjVi08VN242G7MbaciGC/V
0rXlj2D/Isct+zlOke6Go9hNGfT/eWl9Jn/VfF05qPHB67z06rMKvl6WZb0qnqMd
HjjeSNzIUvy0uybJI4cSsJ9NFMWpg2AEYSgT+XktjogOfBDj6tYEm+yAL4jGX8Ft
Z8/fslWtE++b9T5Dpteu8H2HG2jqgCY0zsHIUILfhtLZ4OwLZZ9cbZiSiavW3EHt
OF/HFzkGYqHJ/MWJ0lw6sRptevaiXVWcOvzK+cCgVvQA2W3MM5T3OcvxPmCZuLQM
OyMRFXhxoIEXA5wCgDV5GUMI5e5SgAofVRoOKIdtBzqUDGxNsow1OAcEgP7CsAqd
Uh7Q+w5fRzlkl4FBXAtBwZgPPgs3kfkKG8kdYwMcg9+pS5AsLtxxKqHzvTGO0rBP
t1CK//sKcC30rh17ziLqrb4VqeCNugtQXxrrpOfLq9bWniNF4gUoXvv9LmC3ITgU
qx5YWQN277bi2thr8qK5kNKkFw4OPqq6jx1FW1WGMtFToMUE5w8Xb80g5uBWs80u
77PS5LgKrcme4thHIWXjdW0KDXn/H852t6MtoNtz+kjs3JkuqjYFPIzXMIix84Ej
pfX7Y9lu2JKXlHc1FdWDToeio9IwGAqqoyFFLb2dAPoXZx5dL4OCkBHZfDrpV7+p
fEn2q136qrz73iFnhp/f/s5qbTXfLLirj5cKuSQybAw/JAMzrOzDTF90dbf0fJsu
MJImaqcgMxwRbokQFy2nnp8MPeYzYVBcmLPcEP82jQA5DM54rit5fo/7g9BKK906
91ZiEtI36a0uTElXrjHIesUBofmCKDYrR5ocmuu/LIViv/yaOQycAt41x+gN2drL
u8PBRgxym1meKjwuhq2rBvbapUoIcHUDuaw7s0gHPVj/MLTEjcK4bhcZY3BNQ0cA
0ACgClA0zjGFeYDJfFwXWNjflFDpZ6PDJ2mu/HFMZBr1gD3uFTk07mHE305IcW6A
jyKmGTJCn2pIsoCMiDb88CiHejxEEOOD+lwAW7qz7ZDG7yMRfaqqRk0ex5GyuUkg
a9seoL8od7L6ilQqGRI1paRDcefNhE0V5rvK7Xx8140EkPCzeXRjmeME95PNc+1V
6LQSqvU3kz5l4HODPnqq20KAU8kl4ebXaYohToNL+0lK42bkbRVgsHHVnibwkToz
94o3no/qjp5er1uKOJXE8EVFrqgLYB6OwkkCYfEtopprrvNEBrSgQ+YytyTgCypl
ZZcAud8ZBTE/mLjFH0NOt4x7tZVTi4p2NBI9f43xQMNGQMYfTFY1UzekVb88WtPg
ShRbOf2tPwQ65LJ/AIltMN6d8BEMtE7I6l7DB+32bWRc1SjEoffAYsdTrsx33zW0
vgeoZkNL7oeDxsCUyX0GtlB/QDJh1e0s9bYm/voZYPWxO5b76WsplZpJxMQkt1HU
MRz/1R7lpD5M5Y7XfqCrxKv1hT4Oj77ROo0CjofVFfXbo4/Z8jDp9d5DKHvw8NsI
DWMnjqiLYUiQ5i/LcgFL6nTVBZk611MCmTTSj0YwXz3MKn9iFs6UCUAUQ6qwcN1l
YRKGTyveAhkRH0WBDxzk6xGq7z8Gjjzzs+vh7RKkAW5vlS1+G45s+YIK0ywgjz6Q
9pu4ivNMc3qDERqa8KqHwihT7Qp0CpXYnbfTkocobqRUT9Pp+EV+aiEnKsvYb5VL
Hr/V8NURPI6sRsVAvuUUXOCQakETCvySDLvbNp+QhnpwG0erCR3ZnllAthzQq1LL
vcpSEIIQldfTOHjGm8GBzBcmuvVQaD1J/O4F0p13XNpFj20kYQuJPEm6A+HLPHdV
WBLMqkW2ErlxGB1gmrKaybpK3zlP3ZDr0nWj3obU6ZAl2RqDhRjbr3Bmtb4BMig3
hx8yoQri6IfwY5uK+q0QpRNwRro2tVi0qZ4J5fkjzZ0f5yKMcBEo5MAwgIhN9bZ3
67VZv5XqD0WwMWyNqlHU6eKd8pw/SW/yGGXDlGexFjq8ZOtHoFDZir/6NQL5Y0Px
gT2se4siv4JWP9b1ftmrtri0ji3siIRIuE3xhb9wAWnO7up7H8sMTtqN1GsalWF8
AlLwqAc4uC45nr2uu0UtU46mqvuWdmeDsQFDW2w2LuosJQk08ggRKqhG5rTK1Oa4
n4D/mbu9xG69YDijVMcJTQMlVv6VavGM884BzHDH0+97jfO6gb8Tf2aehnwRnvyT
Z06HW25TJjL7BoHr1rGxSgjlAhsg5DeD0JKGatGqL2c80OC3ckZ0+10XSLmehwij
oquyIuwmOkZ5ISaDM6x4TyfA5qL8/rlVats6UHDxUwOSj1DAW9hZk5ruT9fr6KjC
qLytlhYpABAiBzhZi9RxanolejQ45mhTKZeAIWAdmnR0JI05oPMXF8FAUZq24v8k
9LQx3O9KG8IDwcNgj9wQyH6zmLqcKzMlz0vmUprslR581vgkWn9mxSgAPXbEMyBs
5Y1EOriCdpzCZWKU8Yuk2BGlS19d/9i3B1KFpHYwItOiYwAKyVaHP+Q3ITXhpow3
tKAD+YQ9W1ThztSP1yhLIuqVaCBHwAsX4lTgVva4OLxzSEF0QMa9niF0Q+jbzPAh
AQCSnxZHYB+A2SfySnrprLzupUadlZG3GXoCKQv1k1K2hgoIhX+PKveFL/LnKfTP
jAWpNce7Av00G59dIy31aX1LuT6PJ1gfWG7313s87Yjen9dglhC8HjXodgef1TvF
XbJnq/ry0AEqt5cLCkR/vrn0QMHMdBZJB0Ss9T5Pq5bDcHNW6i6CqSbKRIBjaVbS
jhoLxu5isdht4VHJ9GNiR8uNvNJIXZ3SX4PrG0096kW4augLEEF0neiv2hU73X7+
q1EMp11tExeQyOOp2HM1sKqcdbmujMHJmu8uaKeKPJqZTOWoL8nHFkErEmpA2z5R
llawGlWqMupz7wvdAwFl2btKmjv49C3Q/iODAyg19vymzd1gAfUKT4TwzvYIS/tP
zXpqU/dBA0c+3U2kEka6AROE0QNEViQIFZKtatV08w6g5KBHE9zYthX45iKhHVPC
O/SeuNzHFH1tAockAypDtjnzFIybhnQb60GJvOofRYqlNSD4VFFt7Scr2tprMt3W
+Bi8xsjD5zTPDDQ5JerPFvDXPKMvyh6Qiv7TIB4IfGrB6BjSkl/clJ6+Sekogioi
RVnwenCAlhXiibahijxYY5ZJi8wVeBCr95qF2JzmxBbpjInE3A8q3G8puvy4oX2+
DQUZnl5XEx2WONnPMP6gl+vfbho9M4+CBaex474eHrkdtD7PFPXPwU+Zx5SF1C3T
+mxIuUyuZR1F/ymwL3OKY+J5AUdQI6m5Y18ar+F6ByDWqO43OeF4K7QABbWeLw5F
LDBmk1zffJdr7iKhio+sDfDemEhEOG24INv58fte033sKjmhSB62JFHQU1RmtoXX
Yqr9TVsmyPz87kMyquiTdFDQcJ87LB0GWNQM8AhN9inXP2px/It1ty7+z7M1nWZZ
BUaHSCuuFhBNaDIg6IQs66wTVJ9Gh/ZGkG444oWOIowIHitPAOdcQCFnLg4Ge8sj
7uF/UPH5ixQVLov1iNKnDV+awC5OfXztmnHrify53fBHrrDjtCik1fl1vG/DBZV4
efAsmEZFGPgYuGlRXhZQZlBqjqgmZUa7OnA91/BHY9RZakEzMAS364cSti/5GaDp
b++GhVlIlRS/O1UmxkWvQ7XEDU7yDByHEo3vZrFVCfKcn7SIBTPFbpahOCnQ/NIW
R76sHY4QlcD+/x9vmWO6XiPSPzlxEM7m4qNwShyAjqAow0arLXhZZ3PnczMsJ3pK
ms+nq0sw1s7SkpoJUaEJZTxB7TuDy9nbDkjhEN4nrn4nb6ilFrFi/P0rgIkEt/W+
bbajx3u12zkZdbfV/Nb9GoPDfZROrc+RaMeyzVlPdhtlj31NYslYa8AZC/CLsMbl
bwxSBUxZpI2rfmR47LRS5t8cQTnVEY8ZsCyeWfrTvwxhkRi8wBo7859jiXj+KalM
JTruPfdI90JprqZfF0Sp4y3WRNFtWl9HRr5HbJ0TUYIl5YKde16ovFH4cpLI0j9W
mrzngQBPcXlSNm4vqEdXO7IIKucaGPT5qed3bWnpJKKr+4zW2TFplw/kK3fi0r1I
FGVDl27BppV5xAHVqNde42rKMxx71aa24F7CuoMjAo+C96rIDbO2cWI8pw+6e6TN
ovR3/sZWQpCO9VeDukHW+H1CEdm6pUfU9H1QN3SL31JRX99h4/hmn+9sTqpg9v8/
gePRt0Oq7wc63+Db3NhfyW3cEmkBKGeIxZx8UbIg7V3XeuvX1gk1gCbqBjeUHy91
iq4czOxrbhSkgDlKLARRjqhOWhlCKp0KJeauXdRPaSW5mslXahyHKuhzaDLoMBVH
WjG6YCNR6l18jhA00mR2IuywenIa+qktoPLhtGNuUDhpXG8t7Uyc0JdYfpJ6wZ2e
i/qMDt0Lv64gFOY2juIXByzB1uzN+Qxqv3EYXZbVpL21J058PGV12+PfOzP07jfr
sQL8cqccjfkvO2iZ+0HkNdD0WmwWKgQDmPTWihP1Ryf1BkgjOt/uTZa0MwUGZ1jN
UVF4DTjMtoS/4mohon3INCCIPH9rep/Ed+zXMqWDTQ1/EghkFnEZNjWbN+9R/JPe
H7RrAa6TonTTKamgvyLUY8q8vjJifz9SFx8Z1OVD1Q7xaR1B6lpnwRshhL+8E24H
eUcNQ4Ip5Oyd0zRnTGv13dCzPDN6vJB6AXUoRC3+V3B+n33BIDCxy0nZ4hJOAjpf
UvWiwFFVcYtQemtJda7yc+xMp9Zgr2jhHV/jbPeGDvRt6NJrxuNL7phLs+GmX9Vq
AgXqjVd+E9GSChSx0HdY7dT97E8MMdbhM60Fi2k8N32fHOK+oE6SwGDIN/S2nzxV
5uHKulUCpvGJvVmCZwEr4hMNe30UfTH5rp/D+d7UgE1UYuTORUtgyCtJD7ynSZVQ
CKKm/80vlY50MKgSMrPl8eYMUvF2ApxkoticjDmi+ZBvrqxMJNsfUEo0LIvPUjnj
/503Z8+Vl423MzYDzYx4ngOZT06VP6ILz3N7Edmtu3YMUntEX/2Wcl7dXPirIF+A
HWlYikijpcHHoCjJZCnOQg5uznj31DZnEppnP378UjvGMybEq1FrdIkl0cCi4Rr0
2ZIFi88a+KRmfZ6oBTGDa9yYQXjoB/9GIi6W8ebBaMZ+5shY9btSCxSmySgBdosq
S0WuYnuypDv1iQbe4MNfb2llsZmpmVYfaE87FDhMHwZ7DsTZcmd2RPP+HJJd6HNf
xcs5NYtJcwRggsqJiZR1BOIhRaqlckzD0S0hBxB3EPNyeWFgZ/e61seW6SuMF9a2
TgoTvu+yQD1Ox3I+phXkV7z7h1xbxvfLH7GpF5Nt4T2l4v7H1Es1vl5ZTWm1azBB
MidxOeN4SWpeUIMneF++1gNxMIqTEOVqRUD4lG28N4FKrjuh6zie/AbTTzddTUm7
Jyc5XBEYZe8YdwvLds+LRan2iH3sska6yt4fWfokqp4dqncf1Jc+CLZYb/GjxOlK
rEgbwGyo7IV/43uQG1jHxx23rz95Q1T8YCBWfCWXzx1MICEAsWsHQyt5mnbUevug
diUozxSscTN+I3nPznf8EH5O8QoMtsAhmfM/L/5htRNZtRFm4AhFe5HvrzKHXpL2
lKnJsK+tfE2FZT1S37VjfKI982+oaM0gDQd43yxrhFWT8qu0o2KzbgcjxmUvTXGj
Ne/6V5Si5IisKXtQ9aVn4rmH5C7b0G2Fz1pc7wHiVMb6GHtRUxr2+9N/Kr7SCoF1
5p8cz4vsz09cCFMk2Iaw5ZiqJZxjMdj5cw2/egRX88CHYJlYXtm4B8V3Yq0cBnwc
ls5Q6ghScHziRcy3NWEbYXFafCTKYO+vjSlVQfeQwM59jB+Jq3AIR6oL4qDbvXnD
4KWR3JNtk6+XbfGwWaFozxuYk9qzCJImBKL5nCKJuoxHOvu8F49FedDAYNzT8wNK
QeNpHlf4ZYWMYZC5ZX6gLB2rUIO/9G9cU8FRYZi08/QsMaa1M+SMkjTuJlvqb+p+
GQQWfekMvl8scuWQyuQ8r0fPV6QBDGu2bcFfC0gamFVy1X1vmDd5L11mH522uWWh
opNbSGSebkelF0MZiMz+jqqnSy/GArKX+tlzUkUWqeEpWZ4yL5Y/ZDj7tEkWaj0Q
Kd+R9Bjg6b9xA809XtlwXRM+yr8NhgVfYZyIB9aL0YXOEmd7CUIh1lvVfBkqbLoV
2uLaP4K7IzHUnLYysLDd/x+5KbFumx7Pjoqidpg/jUL9uUgAXtjJwCjvK3llcqIr
/TOayPSkjsh8+l6sV1jSQdbS6AXnpoPmbvDyNUJnSjidJXdYZ1W5zpcuLBG1DsHF
cglB3TVRmvm/Tn8yKS/Gdcg7tTkVHO5GN8IyiCabVek21K9YyXaovV/7TBr9a5ks
4ZtrbIOCQclc/H52gZzqFfsRAgQGjJpJFh85grFZ3QeQgq0bn/dRrmH8RFPRIjbU
NOCXNcIHb489Ov+ZZ2YFWRVl10RqxTrmil4A6wm2ZB+lhsj2bKusQbYE99W9ly+5
v3ZIJ93vJt/y5/QiF4QOpsgu6hDrj7nSJOYDUrcLfkzgk/cMPtYhC0mmns2seOOI
+i+bQ58sar+YyqRa2Fa4HHscAJTo5CXKoD0nGrFxXihh+Jzkr606ZnFT6BdFFqJm
s00A0D1TE71JK9utcPoLEiYwskWEfoeu8aT+NeZUEG7jEAWv7qBbw4B3tvoK9tSI
UN6ZTQdoW5iBOTS8zKjAKys1f/oLEtEAcHk1Zj2PMF/WR4PXkMRf/PO+VzDki/1b
KBD3Zfram152p1adF3rlCl8S1v9Qe1xqYpJbmJQgVUMqZGYy7FwMCH6TsBmDexvw
n64EOnLnvZqBt88tlEDsOZLDXASsl493tjFwqmozqqil9WD0cPbbVNhv0ZXL4Y/Q
iW+BHkTyCsxFO4kU+2VPszD8ScZZDfbJ0tadgXkw4OnZJ+PG56iwjENVpcsAKSew
z0ZCmdNNh3Y/pEyw5zDHZDlC2qgH+shZilSBVD/s3cEQZ0+i17xFMi81vu5FiSeY
2/NcZcu0zaXGbxzuCSiUGF0IVUja68mpPirHG7LVA16BhTZT0bWSObD+TTJEo6cs
Wr/j2ewjIQ5BkWqLK8ddyqItTiJWi8WbkZHiajTh9IEMSaG94+DlpdyNF04VE5gx
DSC1ONtrsqkwdnxS5TK91J5eOEYRtBBk9AdYePTPcOo8F0sok4pco6S5O51h8cUp
LNQwg52EPvcrWBVa2rlnXFFRynATrTtNVhq9IjsuWPgoMixJr7YnMzZAAuoJ5rcs
lr+O92YST6KCSarJ4L4nVn1/kwURXBnyYqR3jSJihqlBC0PSSqmPDFOFy/2Q1Y36
0syissCFdgWFVN3XQHm+BYKdT/pnLIg0Sb/hfvLqAKV9rDhcI0OtcAztvxwGdmgU
D1yVCuG6wIFRJz5kPWnn9KAgwFchTHxPqTKpnWa8SmiWanq2n9UKwUFFw1PxUGet
4iObHhX7PK7pVsuwLB1CjGHW1z0khr3XVzLazmDdTG90f6QRgQs+RmKo5aDnKAOh
O4lE+I7OJmdV35AIwgGcg3J9kW4NluI82pavm4Kx4WyeVoM1CQ3dEI+GAvrKqXZY
gtoeEvXf2AOV4qJpmILI6eey2KurQ8gtL/BQBovbrK+RhCX680HGD2Tk1j1TgSTG
PrGs04vvCFquSESZj8noUuG7NppKRBMYQxYmkdDOUN4oUQV7ObKBMMCEUbRDAcjC
KMTzQIJB2s3XPSaH+3mcUhFMSKilMWu6WAA4izGC7rF2Lp+h5FNhW3wyk7QPEOnF
1i8fYqacCCZH/oVbJaCisxs/GdnihuxthLTOET8pV0aQ6MwOzOn42H4JxBfF8lU9
y4fZigKn0JXRDqy/8img9282vEGxvsJ5VwPrwmJltX39iEwM4otVtV46Qa14SxF8
oy/V8VUhzdzgtP7/KukWYaw4ukKLGo8zYL2Y1W4vCpQxFl3BJRb7pPS4jbfarjjz
UQ666LY+WlnEZ3yoxE89MvCmMO2fSRp5YW2St4r+vQHTV/uv6Q19jJ+98MwvkBbJ
g9L8DT4rUfne/deJ905IlNiRTC8JYey5a4BW513biN1QKRdyF7qA5jI4aRXdZtpw
QFbxMRIcxVxPQNZZJKMb27/LbRuJJKfbkGfNlV/ddnMeeh/j1hus5YUFxCNCEjYc
0vh0MOiRedlh9xDRneCpRKmXnVD73A7u3ZyZn/sz0nFTvsfJyPp2N6U/8B2atWx6
gqhHypY+Y4J/eKARR2OQJ9qCdYfZsSeaEIXYraFuoE5Y4j5g8xfSmtYly+SHf5o9
OJNlZQ7pVFnZYbFppp4VG6tB6Iiwr8B0R2vxjTyhBMcw5Yt8+QqieoE3taCPYu2p
+JDY07YURBrNxh4ltCREU1jI3UgqvPscjijJyd6wqXINIW9qn+d77EVkbLkkObih
xnO3ah9bi176LYXYo9rCmCm2wJEtiACmXf+zlrSPaEFhFAL/kwBHQc4mFWH4Tcv5
vOJIyNGoGoHr1SKc4rS+6YqV+s74Pu7ODES9EmkitO96f/iY0wN/fugvpOUiUA2t
D4EgqFqN1yXAFD/1mbjGv4s8YNWTTQbY+ZVghKq3SHR7GCoUG3IxAlDDMP5oNyAn
iga9+Hw2sN56MbCWB5t3vSxbtrPyjukTTtMYg/30bdvczMsilwqrI6UYCFMTcEGC
83salYzBzkbS8OjcTPMQv3o+UF/5iR5T3gkyLvk8oOPr7TQBfrVQ7glf1J+iyXHj
a7tEs8TD6GsT4W7HwOw9sl5CPecDzEUpim6+BtCES9YgFH/Iqu9Ro9dF8nz2eU9Y
Oq1i/B/tlWwUFfzkqrJf9BrsYhhE6moVx67sZAbsAFrAOPso9zXfTq0RbzOVkixn
1x+KMkRn21PxHIJdvtJEtIdGJkHrH814OvpUfMv2NSvju4NT9HZdKQf3pR0jbDZ6
li5ZwrtXBRLP5Ogqywf963GQtZz2Qdd8S0ZhLM3r80+73TQX2QdVrzgQwHHdDBPj
Icdmsnt8epmjx+yP9EpDp4EpgD641jW/YuOtz7clAfil83KDql2c/QHYkfzq5kr/
44jY+LV0g0SziuhUjBYd8v74NMHjqYjUtDIr8GVqNuQkBA1wD4j1/QCMJp6tods5
F0KgcspPGOnIkCO2f0sQYk0DXsFEHRO7/BbnSrGLCpnB56bTvhOKEOR21tZFUzo/
SBlP8YFaw/t/5QxCUah730g/BqWdTp/n6luSTrJFcYH2byznSWqHAJ7RPe8hvh7o
jJwsWJItncUi/0RUUGfqYGiFLZNHnxiTToPX5n1uKQeR/nT8+WzOx0k0UBsy75yI
uezVIV0RQ+j1g/FljFWQ9O53o8or2ASUL6gKrE4vrKC4u1jxjxIQUyRmFXCekoN8
vjruj7YBO3ce3o4WqcpXNXYfzga24ykb/DXJHtwJbeK0OEyra6PkGtUwsQ1ZMUYq
nSyM1NECNZGhXTbUjmgepUF6jDw/+8IsOW3nqNItz+o8AGk0P7d9yXDNHXsnhuQA
szyH+B8q/izzw0zvJO2Yu9MtrwK7N/m1VFQTpHovQG3dbAVtTtZ3QUpZFbG1oZiD
po1VoXRNX83xjdvadTaZyYAA577ZfGH6sh9cL2kdlDTu2Kd9jze5Q9/XSwdvuFGS
DHFm6kN8mPa/eiqoOm4WD6HbTAZAsEs+Our0XDTUEjzBwmKFrrf1abMObd+5j/S3
LaOyjq48OwC6jJt4g21i+Ka250wwDR4C+xEuoRwqWA7StSuCMbJTFkKPLjQncSFs
MOAe8qjkd/HAGfKT34rI3khm8rlDXtJOKOz2JHM2z0YAsTCaVMn8Zi1u8vxT0t6l
I5CA91IiaYOu1X0hhrlHWkk/d9by6n6Zge7S/+2Cb7UM7AvUrONREbhLSIsoxYEe
qqr88VD+SyY+LNFoaWT5L4mDIVLmApglicvY0ByDwPSvz1Xm7fHUfoT3LyA3xfIc
Cv/Oo5lNkc4A+NQVggoY+i3Lfo5P8rzEr/ArF+USOdeMx2tesWXJbKuINiqRJrPu
OxQk3RP2fsDZ2iXqDatT8fWVaNfpjWSqCOfLM9i8HSh1Q3p1LaHe9gVIIhoQJ5wG
isnfZx70zCWsIpTRPlFk5/+CjiNop2dio1LePGDg8gBpFJ2O0SfnIaqJfHYSgo6p
n7ILxMV+OuWQ69WHoL5KHCVcZl83mVaeIEbrscqpkzQeUWmPvI41WFUydUmglxVy
BWiPyyaTv/yrkbn3X0KU37x+3glSxeZE2aJwuMCtMrA2/t7pMGcW+Z17u/hqpHeu
bDJGeNaZlDeH8MCkmp+qwylw1lvEPXqr30waC9JzJ9iFcW61ML91IrHaTAVzh44u
W6csfBhn/qUGv/HEiEWT4kMrnYEsJKhpVZ+veaoVZ+ypixnTvhyIcenOiOiCClq/
DL3fd1kk3GGpw02Txj/IBuICl5QaEquZEHxLiNyQPwYpKxWZVjl7XeaDQ+0n1hLF
mrF6/rf3meYQ69g6Xohu22btUKxeOVgo6fO6CrEg5+nOJoFMbWEHc7MaGivFhL84
mLGDc0oLiL5TLJvq+UNCTCc0/+BxXn3I9FPj62PZcFZUar67+nMWN1J1mEXSc7Hk
JkC9vZ6ENznblsOckDfZjTcswjBpRRecNOo4h4DAm9RqiH5jKT3sS0TeW3hzWFxU
Zc+AfkceFkV4eHpVk4ZBhmGzZOSTxSYoKzPGrZk2+u1UVr6ki6ljJ4WzmjUEGORM
g3is0x0I7oWfN1/DRokaJ7GUnGKZ6xv5A2PNb5rhZkxKhzXi6Cvq1ErZdEU3uV9E
Dg9sqV/WfuB7d0tqiDhkaTspnnMMk2S8V8m7BwuHkCUmeib5OowiEzXMRce8ayhO
KkFBzVpd1YM+Dm528vkUMwz4Zd87+vpuhT/aX1llz5GhY4Xb0yvx6eomQ0T1G6wn
wXKyfg0Ff580GmcoAuLPBOzal5k8XaL+Mr/YpTliRISnWTXxE9h2Dm4IrPt0iqZo
RZTkJocl1ZBZWn0iBDRg9vkxBFp6YxCbecjsYWMy6RoaLOfv8Qkr1jx4CAZbMNmc
Riomj1edqigLiZDnioMv1yq1DyUsphw6jBpXCmiLdRtOF++DjOBrzzUUQvbuL+Np
GtiBIyxawYubAWNwyYumUDGTjDMHkC57MeK5I+mhCh/UB0mxklZnDN6fMD8hig3A
u5ZKrRH/3H9SA2/B3OFL8IKzTtIngSCKbJSDuStRuI6FU8O4/B63Agfag+9FSjlU
QgLGAJCNf/zhIP6wunHOhyMXqZZie9q9WeQuM2ZISwMxKkMW9Uc5r3CFTg5dhl5j
tlbJs35+fEMlPw8uhlPyyjAgRfxQV3Z6QVLVn5aNUCzxAQqgTc9otMKIrIVCghvJ
jEcF5tAb2LlREIGshna9kuPXMeLzsK4nRff/u3wt59MaQ611qQG+Xstx/HpKwtje
taNH00JEhiVtjeOxab1iNJ6qExGSrG4BPwE9plwoAaxB0GUuQgRhRjsvZ10k3xf7
9m367Ibf+04ca0D9Rq7RRBQszOSw9VoHNIIP7n1foSlL6BWGSnIuN8cU0a+t4nr/
li6iWBMaGTp10FDGF1gcBYtWg87Hx/Qtp8gliy3c74Xh8gEGB0rNhB6/7NxLoruw
R/6yvmBBorKnxG8hCxE3fnCVF/TI3PjygxB3rax+0fGOYg4d1+mBN75x7Fcy7aDv
hVdJPr9Ux0smvG8DxsUV56dBF8KHDENpgl2lEEoKSnI+HkZawIpwt5Osr95gPE4e
DVEPWommw61Fy7bJCNQfl3Z4Pd1YYMA6RUzsYsrb/3XDteY130Ocr93pljcLcx4j
kyjUdNNM4qzdIcuFNHXma8DZLHmyQcKkDy1I/lnoyrWWUnBm2g07Y7x/1oWKrtUs
wRwPpzbjXZWoQS6WOtFxM9u/JtNH4OHJAHCjp6uUtaQ9L/3XjBvZnua13ZkZ9vql
egLPxJqjsk7nfDNk95apyP9SIPrCiFstpAY+IM2JTxugy7OdbcX29iwL9JlTWtHV
PwfvQgpow9S7pI6uMZyuWijJCNms0UEF7H3LK7xgimdyykmwOP7yB8/K4afJo9hT
Rx+PcTPJn6bVBEfrbs/ePnprS7VlgYz9UiTc4Wp4/bbFY7lNJvWHi5HsoJFGUZyX
cMGjcMgh6Nev4ZF+f/lWZzQbU3lp+orgA12AciMhmPc0oAYskkitdqTYalGCMu2Z
s17aplDKUuobfbjUA+lpwBzOh0jDB+W26611baHiykdezB5ab0SLk/ccpMsjNMHN
9Fr6C6khG2pYt2Vo7VFX0cE3AhKCxZMCglw8eJT/S6l9uuBLYsQyzXooBbOHB5WB
lgxoTwMKZtD+XBH+tuRQWtwjO63r/PFqhUK0lktdeExHmNh8VmdNVK7BZZaHxQf4
fOqNlnlz8lVDQAg8An1zsIof2CRO/p75wcriHZctx1JPSe4+Egqm0AelYA/4JRoB
pMSSy2VrRVQzGUqAtJ7Vm/FQ2WXQjhmFXTvtCLqhINkL5oc5QW2KSRDnD7RKLGIL
wbcVRGcwWt6oi+PnWfu9o9D8SzKMLVIQaSgbpHYX+QQztL5yy8BLaVj2zcHrgLjW
jD1fMZBVdXOhtxIDymyIz8PfaWuaX1IIozYcS9icrdLTU10MxDijyRPm0rtM4oLR
lFzG5I8d59NSCs3LZx5OKASILcrxQvRgGMbF6h5p4PHUZ4k76blqiyUOFrIUUowb
b33bkbE4XXY8mfr3daNYbKF0kF9TaChxWfHHDMvW4KkN9eRmmUmcos4NbRPpeyGE
mAH733jseOvVTU8fIQxRbpRrTE2ROik13EzJhRlbCKNw08JLHB0YvMu7SbCh1faA
Eh1xncH9dvslOSZLW8vdvgFXSNj5NjHg0jtd3+Qy15tXTXCy6byH+gQg4NPJ/BZO
bXMEKRRyQSubm4519SfV6QJIO0JrPDhd3sTAHn8WgcaFkcV+hKF3/0TrlxzPKjEM
zqO6U/Z72XgE3ujScCFxv5YYsiDAdBtUUUO1fdiD2IDYL2y4VGtEcbP7sxfGBLRF
3nOf3bnwsQ09w0eIXLterUt/gtXsf8uTWv5Bn2e6615LkrxRoy4FkB5X2TTAYb7w
SczsSIPpsojYRS73x6NLFAxcJKtWbbMtfemNz94xZ8AW5LZhCYB00FqPGjA42J6d
6GbZEmKuKhFBFK4t7rZOc1SSCDVu1hnaxcGP3vgfLfsFWvQstwN9fYOTNMy34+ta
mIrbhQjBuGW5J1fT0vCw+uUgN9e7M7x4yYpzVmPXy9Wndpq2vPo0EDOeKCjBzegi
p3JdDb3H2hockPwXFN6i1algT1P2B5XZGYi7217KEIBZUKZaRuCyGuPavGB/djJG
6YXMgDJt3882ggJi/Iav6YHaFAWDe6ORqQ7VhQhJ055JicwRXqKLEplGMVRXBd4E
uRQdiP3flvFF+1vRFm/gM96CwJxssJwPTA5HO4kMaYUvRHV4XjgsRZSQyprXLGsT
Lin6kkE8dYueEAFJDLh9RMLq72zNoakCyNmYGC30v7J3xS9RQtPKW/xASPTyAmMj
pajtZpTbUnG2UqsJUlCwKp/57Yv0ZkFquk89b6B07/CkHcaaBXBhUKle28qfYof1
z9CPEqfmUMJEZNTCVaQ83Y56uALL8JNUj3LK0ZHFt7BO2cNv+nfKJiB2WyYHnAHN
XYEEV0vvXVqpAd/Z8TXZcXi8QZ+bS1aSGTLGlUi9Zl9jqRWy2+uyrcpCToRG7yYT
DO1BGeoTqGrmAU/64VxFNjfN0neoKStrRlN6I26BMvZl9bo57yD/guf+altINHJM
P8o5St9qEpBODm4v50UfBUEIDognxnx0IzX/Ioky+FZySsk5WEz2luIL234lbFr4
mkV+Ww6D9os4euIbiIRI/lO3Vakk43a27TI2anFhHBEcKJ6ZS3Nc2GpkXOP6sM3h
7Ts5l9Narv9usRl6zVlRBJMfz/b6QB0oAcf8E+EEBofWq0NH1aTy+fqc+64B+gSZ
zMg9XKPe0NCEsERa23BF2vwJW2t63aamq0KgaUCoT1taz3Saw15zm248pIZ3j0oZ
sIgvEcN1gXIdGKXy7SwfRHB4xpBH7a4bYXMtHJ4uOAYF8VbUzxIaUHTH6vhUDPGz
DG2Xh7FIaM5E6lzbFFDU2hNUBMcDKuii3GCQkrgDJaN1L+baEDeXOwWKN/7EF4up
O8AzHMxV45XY04e/w+R4Isuu6pA3lNqmso47tWNv1QJafBS6//pmjE0yWe6H3O6m
XPfnmWMDRTYUZXCR4SvA+Bg5YM4ThRMzb+DpR2euXVtqqwtIf8TDviHkOdL/HDJN
+1dFckEIIS1sMZKtzXC0jf6BejsBKCjJM2OhbyrMt71yrpa9+zAmp+ouL8UiX3Ki
m+XvW3R3sy4asLuyTjithhIeyBwVuOne2h8scVSOjDLLNzB+fSBzALlLcIGnvlEc
pshq91OjysZPgMl4Kuh+1CHh9QyAB+04aWMXSlM8XoJWFJDiTh3bPh360/ORFJtq
4FBkweR7f+JN19V+PRONYS0+5r02bxE93U3jTHwihTYz7ufhale9edMdi6dG+eIm
MNmntE72oRj1eWdYN5UeDwqwHX6+KdB2BDMhDpDOcEU56VxCTn9/KghJKFgTKm37
bOzw/YZl87sICft2VYo/sDlC8bXemwIax3tYlQB+AjcJ3DzOc8wx0xWZ8oUtsOMe
Otpu4D1/KtFlPMpt0TzS/kplPMA3VwpSUgmgpVUNbmHXPjeXElTHoCf89m58AjJy
JWQkMR++J5to/Tg7IYOLy1wgjNh8TazXfQEUqZBqP8QjazCR3pBZseMmIHD03n3a
Nvpkfb2tJj6Je46e9FyKzKYhKKuJJWU4t4NDOGLJkCVKvYKC8HPJwniagEvnq7Cs
tPc91ddKSdBt1d5iBMjh7LDIOemc+EJ+DDIDZLes4AJ2aXhFoTbZcV8B4ByYVA+a
OB328/C+y2B0UthalbgL5WLPS2j9ZTp4/fZJa6xa6iEfgZ737kj2RjUJX5TtpK4T
qvPfpQLE+Tjh/KqCyfFEKfAm2Yq1MzXjOXDovSPXRHzNzYAyV/MtxJjg6tdxWSUZ
v1F/72KeG9K5qOTtyxPruNG13nRJYYM1gC3G3ogYxBIDhNgvxC2hv0MfHDwHZOJW
bFjw16JZeZjXXfpyVUOJOBcs8W2YCO7LY9z54RIFHk9IEW1T8UA5qDMQwaDlfs2L
BbFLwnfQgZE51Bjg+vEg/8AEGF0Y6icDS7fTjgasgrxva1IieYURJbeiJwwh3L3m
lDOlmMom2YSx3ya0t73VVwcsn6JN2yzzwY6b3zbxHIxcRTHskV52y9CZQPEDLXST
EXap+38scgeTSH7n70Op7dXjxpbAu08yOm7CWYDfupo2NHtz2Q1Pc0ayb/VNR1R7
U/8V1S7S/urcvur59jEbm+2ikSBxIgRPXmo/qkminPHPVA5lgq1vVKIrf71UAvUv
N2HiETxwhJBpKzFFLqvqlZjmv8GWZyVw2NdLDuIV5uxCeMu24dGYZNl9OAjGa6L1
2AgOWyX3nqSfXmEBnFBGIByrQ38hJ2kbGLWPiVRPvkME2Ynv5A8H//vZSED+mDJB
nnAjGjU0DDxMXbPEWTBpikb71P5Bs//d2KpbNuKq0gnbRkNtz6/t1xOqJtAqaHy1
FpaK4jNHWIOT7bAqC+rslWnuvMYxdEOkVMNwAxQcSG3RX08fmXBX98j1MN+ojFxM
K9nsXz1fhDfmAeCs/X6/fuxem7EtkjhzE8fLM+nl0J7Z1V1vQxffppWKnBJczZBW
TY8q6mMo9tP0P0dsqDT5W+jBKwozE94DBBUuzjEDMsCKAGa4QDzyjDAVIaRd1Q+8
6WhTfYd14XaZ7VB97z4TcGluDc9EIdtfzcdSBFI/t70olBWklyXZIS1XwNvJYwdF
xxPk6V5dojLO55aAYzHylc3cyVk/qvvQf14tqmRH6Uj86uheEg+MsJ2pAbi/uf68
l3t37OjGQFNNopL/lShZN+r/wgxPEYiEuK3jYtkpOZ9t0AxYDH5vqXthoN8zb7Bi
pjoZqEeH9uKClC/nSk7A1vo7VhcHifVcHkyCgG4KTFmfcskjRvPTu3mpvmgXg6hp
f9MSrpP5EUQSOvCZblxRrbfjSSMiuOSTYK9LEFY7L7JVvsHkw/k4RXpVWPUW5AAG
rjCkw3hB8KGYKLQUGYiS1lpOUnLfvPDhEu/gbeF93sxJkIBkarvdmM4tNo1A1cDg
ZtjopEDnkaulwss/R7tgTvUN9AQV2F/CEoN8xfdCdo8DJQqeanWsjB9y+tT541pW
oaEeLCw6DAGJLZc9hQl2H3MmaikAj17ixNRLwR2TqpgEBNuqc/aqQAamLMKpR9Aj
`pragma protect end_protected
