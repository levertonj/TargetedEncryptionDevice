//////////////////////////////////////////////////////////////////////
////                                                              ////
////  eth_avalon_bd_ram.v                                         ////
////                                                              ////
////  This file is a patch used in conjunction with the           ////
////  Ethernet IP core project.                                   ////
////  http://www.opencores.org/projects/ethmac/                   ////
////                                                              ////
////  Author(s):                                                  ////
////      - Jakob Jones (jrjonsie@gmail.com)                      ////
////                                                              ////
////  All additional information is available in the Readme.txt   ////
////  file.                                                       ////
////                                                              ////
//////////////////////////////////////////////////////////////////////
module eth_avalon_bd_ram #( parameter   DEPTH=128   ) (
    input                           clock,
    //port A
    input                           wren_a,
    input       [clogb2(DEPTH-1):0] address_a,
    input       [31:0]              data_a,
    output  reg [31:0]              q_a,
    //port B
    input                           wren_b,
    input       [clogb2(DEPTH-1):0] address_b,
    input       [31:0]              data_b,
    output  reg [31:0]              q_b
    );

`include "eth_avalon_functions.v"

reg     [31:0]  ram[DEPTH-1:0] /* synthesis ramstyle = "no_rw_check" */;

always @(posedge clock) begin
    if(wren_a)  ram[address_a]  <= data_a;
                q_a             <= ram[address_a];
end

always @(posedge clock) begin
    if(wren_b)  ram[address_b]  <= data_b;
                q_b             <= ram[address_b];
end



//altsyncram  altsyncram_component (
//    .wren_a         (wren_a     ),
//    .clock0         (clock      ),
//    .wren_b         (wren_b     ),
//    .address_a      (address_a  ),
//    .address_b      (address_b  ),
//    .data_a         (data_a     ),
//    .data_b         (data_b     ),
//    .q_a            (q_a        ),
//    .q_b            (q_b        ),
//    .aclr0          (1'b0       ),
//    .aclr1          (1'b0       ),
//    .addressstall_a (1'b0       ),
//    .addressstall_b (1'b0       ),
//    .byteena_a      (1'b1       ),
//    .byteena_b      (1'b1       ),
//    .clock1         (1'b1       ),
//    .clocken0       (1'b1       ),
//    .clocken1       (1'b1       ),
//    .clocken2       (1'b1       ),
//    .clocken3       (1'b1       ),
//    .eccstatus      (           ),
//    .rden_a         (1'b1       ),
//    .rden_b         (1'b1       )
//);
//
//    defparam
//        altsyncram_component.address_reg_b = "CLOCK0",
//        altsyncram_component.clock_enable_input_a = "BYPASS",
//        altsyncram_component.clock_enable_input_b = "BYPASS",
//        altsyncram_component.clock_enable_output_a = "BYPASS",
//        altsyncram_component.clock_enable_output_b = "BYPASS",
//        altsyncram_component.indata_reg_b = "CLOCK0",
//        altsyncram_component.intended_device_family = "Cyclone II",
//        altsyncram_component.lpm_type = "altsyncram",
//        altsyncram_component.numwords_a = DEPTH,
//        altsyncram_component.numwords_b = DEPTH,
//        altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
//        altsyncram_component.outdata_aclr_a = "NONE",
//        altsyncram_component.outdata_aclr_b = "NONE",
//        altsyncram_component.outdata_reg_a = "UNREGISTERED",
//        altsyncram_component.outdata_reg_b = "UNREGISTERED",
//        altsyncram_component.power_up_uninitialized = "FALSE",
//        altsyncram_component.read_during_write_mode_mixed_ports = "DONT_CARE",
//        altsyncram_component.widthad_a = clogb2(DEPTH-1),
//        altsyncram_component.widthad_b = clogb2(DEPTH-1),
//        altsyncram_component.width_a = 32,
//        altsyncram_component.width_b = 32,
//        altsyncram_component.width_byteena_a = 1,
//        altsyncram_component.width_byteena_b = 1,
//        altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0";
//
//
endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
// Retrieval info: PRIVATE: ADDRESSSTALL_B NUMERIC "0"
// Retrieval info: PRIVATE: BYTEENA_ACLR_A NUMERIC "0"
// Retrieval info: PRIVATE: BYTEENA_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_ENABLE_A NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_ENABLE_B NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
// Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_B NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_B NUMERIC "0"
// Retrieval info: PRIVATE: CLRdata NUMERIC "0"
// Retrieval info: PRIVATE: CLRq NUMERIC "0"
// Retrieval info: PRIVATE: CLRrdaddress NUMERIC "0"
// Retrieval info: PRIVATE: CLRrren NUMERIC "0"
// Retrieval info: PRIVATE: CLRwraddress NUMERIC "0"
// Retrieval info: PRIVATE: CLRwren NUMERIC "0"
// Retrieval info: PRIVATE: Clock NUMERIC "0"
// Retrieval info: PRIVATE: Clock_A NUMERIC "0"
// Retrieval info: PRIVATE: Clock_B NUMERIC "0"
// Retrieval info: PRIVATE: ECC NUMERIC "0"
// Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
// Retrieval info: PRIVATE: INDATA_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: INDATA_REG_B NUMERIC "1"
// Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
// Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
// Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
// Retrieval info: PRIVATE: MEMSIZE NUMERIC "4096"
// Retrieval info: PRIVATE: MEM_IN_BITS NUMERIC "0"
// Retrieval info: PRIVATE: MIFfilename STRING ""
// Retrieval info: PRIVATE: OPERATION_MODE NUMERIC "3"
// Retrieval info: PRIVATE: OUTDATA_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: OUTDATA_REG_B NUMERIC "0"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_MIXED_PORTS NUMERIC "2"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_B NUMERIC "3"
// Retrieval info: PRIVATE: REGdata NUMERIC "1"
// Retrieval info: PRIVATE: REGq NUMERIC "0"
// Retrieval info: PRIVATE: REGrdaddress NUMERIC "0"
// Retrieval info: PRIVATE: REGrren NUMERIC "0"
// Retrieval info: PRIVATE: REGwraddress NUMERIC "1"
// Retrieval info: PRIVATE: REGwren NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USE_DIFF_CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: UseDPRAM NUMERIC "1"
// Retrieval info: PRIVATE: VarWidth NUMERIC "0"
// Retrieval info: PRIVATE: WIDTH_READ_A NUMERIC "32"
// Retrieval info: PRIVATE: WIDTH_READ_B NUMERIC "32"
// Retrieval info: PRIVATE: WIDTH_WRITE_A NUMERIC "32"
// Retrieval info: PRIVATE: WIDTH_WRITE_B NUMERIC "32"
// Retrieval info: PRIVATE: WRADDR_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: WRADDR_REG_B NUMERIC "1"
// Retrieval info: PRIVATE: WRCTRL_ACLR_B NUMERIC "0"
// Retrieval info: PRIVATE: enable NUMERIC "0"
// Retrieval info: PRIVATE: rden NUMERIC "0"
// Retrieval info: CONSTANT: ADDRESS_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_B STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_B STRING "BYPASS"
// Retrieval info: CONSTANT: INDATA_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
// Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "128"
// Retrieval info: CONSTANT: NUMWORDS_B NUMERIC "128"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "BIDIR_DUAL_PORT"
// Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
// Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "NONE"
// Retrieval info: CONSTANT: OUTDATA_REG_A STRING "UNREGISTERED"
// Retrieval info: CONSTANT: OUTDATA_REG_B STRING "UNREGISTERED"
// Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
// Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_MIXED_PORTS STRING "DONT_CARE"
// Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "7"
// Retrieval info: CONSTANT: WIDTHAD_B NUMERIC "7"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "32"
// Retrieval info: CONSTANT: WIDTH_B NUMERIC "32"
// Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH_BYTEENA_B NUMERIC "1"
// Retrieval info: CONSTANT: WRCONTROL_WRADDRESS_REG_B STRING "CLOCK0"
// Retrieval info: USED_PORT: address_a 0 0 7 0 INPUT NODEFVAL address_a[6..0]
// Retrieval info: USED_PORT: address_b 0 0 7 0 INPUT NODEFVAL address_b[6..0]
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: data_a 0 0 32 0 INPUT NODEFVAL data_a[31..0]
// Retrieval info: USED_PORT: data_b 0 0 32 0 INPUT NODEFVAL data_b[31..0]
// Retrieval info: USED_PORT: q_a 0 0 32 0 OUTPUT NODEFVAL q_a[31..0]
// Retrieval info: USED_PORT: q_b 0 0 32 0 OUTPUT NODEFVAL q_b[31..0]
// Retrieval info: USED_PORT: wren_a 0 0 0 0 INPUT VCC wren_a
// Retrieval info: USED_PORT: wren_b 0 0 0 0 INPUT VCC wren_b
// Retrieval info: CONNECT: @data_a 0 0 32 0 data_a 0 0 32 0
// Retrieval info: CONNECT: @wren_a 0 0 0 0 wren_a 0 0 0 0
// Retrieval info: CONNECT: q_a 0 0 32 0 @q_a 0 0 32 0
// Retrieval info: CONNECT: q_b 0 0 32 0 @q_b 0 0 32 0
// Retrieval info: CONNECT: @address_a 0 0 7 0 address_a 0 0 7 0
// Retrieval info: CONNECT: @data_b 0 0 32 0 data_b 0 0 32 0
// Retrieval info: CONNECT: @address_b 0 0 7 0 address_b 0 0 7 0
// Retrieval info: CONNECT: @wren_b 0 0 0 0 wren_b 0 0 0 0
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram_bb.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram_waveforms.html FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL eth_avalon_bd_ram_wave*.jpg FALSE
// Retrieval info: LIB_FILE: altera_mf
