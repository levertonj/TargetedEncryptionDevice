// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
fpZGnzEOOTfzXk8zzNO1O1EOvYKPpdpdrvNnf30AB+tcdicIEC/D/meiOD6T7stR2Q9ob/OHuvnr
StwMLXo2Uc7K8n49gVNfsYUdscQh9+GMlNplFsPAYiNQGIYMBdgmV9JScU0+hKRhXK3Zupxz3rtJ
UR4cOriW9onEOYAbXvO5oD3zJAGxDakbqkXUT7NN96Bk0SzOvb29zlQJKqwZJZFKhH7pauOXn/Kc
6BS5s5GMZZ6DX5Ma9txxYPSwJm8h+49oU/yjP6pZnqXoyRbV8Hy3RSH85Qh5IzcEVj4kDIZlnJmt
2goIWK4L0NvbjcT8F2G50CZhCn4wNxtZGJF1YA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
f6aN75VT/MuBEN/6fhlxwLMtfBsNI2e29rse9blY1eQ21qTh6jhwtlU2+C089SDIPyKgdC0Gy1fJ
Gj8TzfKHkNZmuOtXhaLdfxdxdYAYHAveuClevxXT1kpkbAd+mCGBkR2L69GOZcANME5NkeHSmYQj
UgdwrU21ENTYSzE/0Jt5iQvu8s/lzgpVVkvsQDPjozKpLzMtrJaPpzx4vKoNwJyrCZfvuWpUQLXw
bW+OhIjVcDkQ5UqubvWgIJM4wr78tQ3Y7w2/ixiiBtdENHWENKtMpowWyItarH8vg4f93+HaISVH
+uaOn/qS+usTvZksCIMIDPfvqczDVlpbrTOHt/Q6asq/LB2YUA2yL6KfshIN7+F+QsQlZhKfHQ4t
65Q7wNyEycW2Y2zeSQOTFBreTkRBnY16jA9/RLbVS0R96YBdX8UTndDUpvhW/vg0U+aiZhInn7ns
QVTlAck/ysJEPPrOLXeERRqgHCZszRlNAWDpwUveKgojzCERvlzopmgunncrcukeq8hvw/JjOuJq
uTBzt917PLLmXn0Big6K1YPhzLmRDSmrKRXGXmAq6gApXcTQklLgTn5ZFip+NQAvmoNqZZ8af04w
/qLAi35tZ3SYQNJYPB9F2a6VdcoLFne8yCdruWWnte3cL+Do3YEte4Og3cqQV7Td+ppk1u3Wv9eb
pATL7PXQRWhS+fylRxJQKGcsgOPvxGbqRoOUxjRDBPUkynUWlxmyPXdgxexxi2oM9F32XnGbLjpF
do/ZxNJjhTJsWFXCWkqgtBArXtT7KEA/SnqMHVK5nQiqxebG6fqv3nvlN9ExDYxLDl1C3vv2od2l
h5NR/I36rEabIMSqNPBgsjapT71WvpTgNAZFykj5oO9PbodY7Rw8ZkzpR4VJf2zHOrXUkSj+zQ2T
PH6RsRx0R48iCDe5XsTPcVZCvMSebekciAZ6yRgShLaJb0eaevNlpbDyMAknr5La0A3UiFUKB25E
zfLA0FpFPHBbzyF8xXEXEGXfnNCbN7Hhpb5bQG7oN9xuYBu1/nkvOW1bfa5CMXf+4FYU3YJH13b9
TIyY+YKIsYPMqwitnt/a5A1dDMcMPiZ8KKq3QbvlrHKaJWXlurw52vomVYNHhhtkyD203zPxx2EA
ZnkQyGnzgl3G1Ox26Kbv4LQzHeUcyzlxtgx+4VoJBL7mr4OsUmJ6ddUvq+14dnWKzPW36oEtdytR
M1OIQaMg+duPcjn9YW8kPyS5xjWFaBoXqh0RfUOUZ6q3YPqD9T17QfdWfWmsKrUCu3oAyoBeW1Js
Ckpqu6mtqQ0LzxvPSmsmFEVw8iRce2dW4OJdptzppHPT3wg527kQJTp/r8VVv+KY7qBtKiJLPl/G
g1QvcE/Kx+L4+gMqHklnkbfPbTm1OXJxoYcdL4PSCqaA6tmfgS7G8C7yilliIC8tYoWLAdploSYK
xkLXtVnZRYKa5NigBmNilUlGIROO7b0IE8A7AYgRDZmFu9Nhcgk/iiRssQrqC/BEHQZaA7fkQ8L2
BI81Cn3kM4Pz0mr/pEdzSBaTc/7YSz9kjmnMX0KHenH4doIb0bAfPlPasAeivHIUSqugx7Z0X+lL
rqvJiZLXlkQDsw6F5VaI7TsvJ3gH8qfcyY0DbhGoGu4iQdqraTyb0bTK7hbrsYbIFNVCMBX2L4Tj
XCA/PlPw1ItuxpaaxojaIO1a+VBPJ8q8Sctx+9hyBIS8ee5CqOj1SKNN/hAuwKktpWyHZnvQEZvA
h8TwrelXHDju3if7GJvkcl0DKbcg72kIKKlMcDZ6BWZvEdnpJUcgzDifwHCxfjJItcdfXFRxrxfQ
vRDZCna4n1Rx/8JyCGtPmsqWTv/AbggdjZVcpcGR9kqPe4GPf9qitKBy8RKwJ8HhR3mOuUGPxc4B
+wKevBUK8uxH0JhYoa3r3P74vpBz4lvbhi2JpjNGAp7Wd1EdwuqiGAPZypo2zAUYOFBtdklENQCh
xdmv4nfK3Hjmn1WQMJJ987WetEI1giC+5rqq/sb6vId0IYPWxLBazqBERiKFVJ8qv3OUksjxWKf/
wBaO+wKo1PMPsMani40rdSgP2iTJH/P0eQykcUoNd7Lzr3rPuzVwgG0Ev78ykiiXt2fwzpvf5Evr
I3eaRRxbdy4g68/a7jZJExOvlx9/gtDz6U2KxF63O+DyLVHlHVXCF5Vb1Q3HJE4L6JoiFDaumulW
8szssdGlcW63jv5Yq+pKKFdAP1u74+tpNG5aB57PX4hQ+YiMP/TLDMncljlxxFSrZgJ8O/LI558W
6jnXhjdc/og4BT4MCBCRs0k5l7wQDmOg6PBTJkcHA0iSwF1bmVCVnsi9GApMuk1HIZ7aRmt6FLFs
TXTa5AYRP92HgZpk0W41YLk4Wc0M+mqKEbMJb1SR1Hng/pi5RJPKm1ZztAbCDqiNxDb9IR+udzk7
Ix3httg0MM09raMlxPLOQOOjHEo1xj3kd0x+NlGkd7QJkL3rwcx71mHen/g5C6N7Iqey8QhW7ooP
FE4Ybw3IAxibIvTvrUg1sYjQO7yssfGTwraFxx++MeXPn9SRvtKGau2pR7kOhI8ZNdouTLGC9cuH
16uvauFaRfGQI5Fd0Lrh9+1K6xQU4NhOKuJbmFvQxBnCNMKF06WHFpHvCknmRfFkpYBJhBtwx3+v
5gRivZ2XOI+mQhgHpKsRA+EQEEUuEKlbCyJQH5wAVDb4TtRqyTRLZScFW2BwfaPIU/uByk03uW7N
Rl9KMyv9bBJweRHs0o4Z7Df+FnFMaeRDbHRXhGL/t4lYbfzpHLDjRsDuHwn1y+Zu2DPaPqMjmaGW
Pl3MiRO6FBoOGp3znx5wmJ8bPTWOwMZ+dX6no2Q1KKl7wJkYxeOSmj6H8EASQQyddPHyMicVdhHf
P+001NMs8msBqfKcfXRWywTTlVdejCKUQG9lw9MMoD5UqZ2tIEQqvP3cXfjkkvn+mEkLwu2GSiJL
75oZQ6eiQkicRuGvRM7D9AAICS+VCDyWi0XMekw8IJbSrkI5c6CvFtHFUvUwJ1mlcJDDz1ydqXhl
MkTKLU/yhGpPxSKXzaZfxe87cvippJRIBgIuP+WT3eof18yzPIuWeP3yrHMlUSq8InSP1d69ISqr
956EmRhx2NXwXEKD9xtDdgYRI5CPC+u4WXoDojosDmvncayMorVvmTyiefzfyUjgerz12cuB9BGW
F/jUk26wVwo6IDcWlgFHXzFuH6tGvWNViu+1DVG7jiV6WLpC/vpArAECCheHJ4MPcsil/6RoQtbl
+ipirtm1ICpkH9ZayldIrG3X84tredy9bLnk+0/AfBsp42PAlyvz+dxvfFJBMB4wMWwM9hKoq5KG
sh+NYLB3Z2kHZ0UcytKHecRBV0r6Ze0J/nk99UxAvzjYFt8nf8L/iJFoJMd69aWBTsmuhZ4SdzBS
2xWERRUM+H7BXz3fahOfdDGICLWoyKY8QkQLqickkPnF79tp6SHKXRxTxvYR2EoMxVzVk/VqrRuh
x9QYDrOu1jPO/a/vDAuST1iiNrLI2ZrwNi0+I0YAn0Yj9S5YNjbiSDq/vY+dtz89JTbV9FuXUSOh
FUgvvl5BS/GDlm9D02w9qw9gzjtjMxMnUdd7z/UvRh92H0z2yWnEabjq4HAs8LvYigacVQIZlnuZ
pGbwolca+srOfoqJJuSGXwmieuOV4hI5RicOTiGjZlT0x5wUBm6m0QQ6TSIZUpwHdLugFooDQT2O
AjWgR5xWe2CvK0D5uWJym8+zQp0IO6Fj+Ep5ujLWr2pZdKPruX9kq5WuPa/2k6sW8alGwD2yY/MH
KW6PGL5LRMH3P/gEDCpgtX+q9wq1wGUF1sWAH24zJkncoB2K8DLDTb3SXVy7HoEseihojaOu0f5Z
fu1OpV0I/BQMfpIDff0WJriZbMT/8kEZZ79cdfZhT8nXBFg0Uu4NrH+cj6orE7GVJX8MAJMCQ8oe
IBO1XPF7+ovqqW95n/yks4nF/c1oSVwHM+VHEMCVjA5XvuBRE6Mnx41zu40UJKdceU74tF6LOErm
MN0rJq3E7swFlE77vkiZjZ7H4TDk2VWH6xVkKgbCXUeJBiH5S6kEVpTS7cmOmH7LsUZRKZ97Hng1
dKY2CfDBoDWO27jgf2Kz+aSv3j7Z/JDLtrQCKkIqX+MD6IJTsUALsYlx6lheIStIoJdHv//DGmln
hol8CjKbhmLobN1PCdoPTatQW8HBOcBFZ2fKcldGCeqeJxnM08HaimQWNpHgrA0GQGjAUf3bh2W1
o8EhT9B/lrkynVnpJI85XWrwRotwoEWbIHVCM5A5j0pp1nOGd8aYvDJOmlbyhxpDVPx7kr8upumC
IgY37sWdlbTtjTEs3oGU8oEr0d+13IHNWqnObOW5lG8lc4HzeLSbPltBdIl7LCr7IBEkmgKJfWw6
k9xglRH517ZCbrlsNIfco/A1IfYx5JBRV0Mx6AJRmmg2CCvR+0M+/KnN4rwJPyrlkUZ181L18kky
LJg2EDkgBFA1CuMCho/y/6qqyIyyPmLIj7YGlDsiZFQFLDR/tAB4RW8ueIxx/ePSUzFw2OD2BX/X
bZJPbjvjVerchnDZtnAOj6w8OucPXHu+vPqrSvDhJWHnLOaPfYkDEI0dNROSLHXw8kpMG+jqdvyo
5WZkn5qco50KVBBWhIGb8tUlKIlXdXHJof3D8Qx3JLZYpCoidUA/XNxewM4U+18bQ9m2kgQ18XPe
WrzA1CvgHZdtA4fG0CJycp8wkctUgxkxqJmVCSLaehcWErTv0/jLn6aSKLafr6BzUNpvLFf6NyY8
3eIism5J8XPnkpMj+OlSoAjztnKGVxR/eWDQXKQ/m2dJtm7728hPrBwb+54ASGUkU+cb8T3VLCcp
ZZJ+XWeq3x0xVnv+mFkuhuoViqFGOk3i4YEu+P3AUH/GtK+kpnQJJvqXqhUNefdxIzBebuYy+hiE
hj0tQRsSP4WyniZ+v8PnYla2KlbK6I7IIvrMk2OBhLG2dYqwF3cqTT/G6je6PkF3aWjSz8vmCs2Y
UzWAiEtJV4c2OWW4k4a4jwPGYetNUyDPN3gjgG+Fjr5n5z/Vj8AHbCuFznEOsIbtUdmtcRsVKh1i
qJCcwlEqksTARnIlk6lk71SYITAd8Y8I8OwTk54lu4o+2SFXsH0fWHFk5u1CelTYPdN0FP+V3a/Q
eIKR9kXBPpn1/o2Hn8N0pICAWWYPlQr2Xsl5Y+iz+Ksu6A8R/XNVHjhUGJDoJfBPaUWDcOGop+l8
va/zPGQGVnqjBGBhiourVsrpkBXZGGl863jq2nw0CeEOwNpJMFZul5RWl+oROlP8L8o9YUFMy37q
zOYkAR9G8SRcFG2+HfQKJ+A2R87vE6FWTEjHUmgA54NrmiHUbn2O/tgWXDDx+d8OJ8XLx1MTYlNs
ijkEq8ftXJZ6XGASapM9wsOvygJgjGv/7pv1os3t4bnyJmW7mw0w3xDlvSDvKMT+GmH+Z0/xyfPu
0hC8EuUzSU+D6Kt9ZnVebuqccQoghCC32KncnJTeqpnOenNhgRPYJpBUmHwhiOeXIbCOaJBjce4t
yYCky6u3ZTO4z2XEFsAEib18KesemhQROaVXpGaj3F2AtPme7C0D4PGganwP0SBdbV+FowKPn4Km
7fSp3Eaf7GXe5532gHnTvhFXpJGJo9JD+dhU/RrrB7mIbrih3e+0xmBMcsGfX7OXhVPaPrIrSGYk
agfTQUbOMtfbeo1qDvD6x6NOn7ysV8KKDDyhIpoj0GT8L75ci4+6tJ8ISIe2XfS2z4VrjPENYDyv
Za/f+A0mbbX4IM1BBXGwh8XONVlsihWOKEdBoy9IcDkEF4HObghpzHwlWQO/zQQ3VajLKcJfp2Pw
NxaNxp5l5BvovY6T3sF7nd0KkRifJjG0oy5DhuxXmQCJd595GmfUWhB1+XGQw8ZHqvm2lvslNexK
/SuIEANNiMsvyHjaG2qGXynY9bbogde3OOnAkhuieivfhhsitcfbV0R4L/LyOXlBN83/NV58tDHx
nGSqsc6ylBNMziWwHsACxMleijIe5j8FhJWXVu9xc1OJRaTSR+cCL9gO9uzW1xMYf74XnWnwRWLL
/KxR7jxebXCUzlwnP9H7f8hLJ9I5qJkSHP1Cle1jM8Y03z4/eF+FFQnO0TuxjrkRBp1PQZ7Nt3V6
FR11ebl4SalmCUw7GPny4awoyLXEuIux8jTXe7kpQXpfH79hdvMMDvTNVKhaSmb5x2lmEmDcy3WB
2IAMovDfl3Aoveos+kiI+cqNu9COt0CQW5+Mb9PMO+vbs2zUr7k16B21Mioc7o+5R2ifVq7bVGo5
rbvbel1htBOOdZ2CVsaDqilf7FEtzDo0kS1FrNHwmJGvVBLtRRRJrFLeQPZS2HVI5a4URZhQOoHV
aHwsDI5Mh6aBfotRmYCD0gCUmKkOb2QY+bgv3Bo4NP5+MV49K/MzVYZpxK58h61y6pW7apCwhXx8
b9W9JwVqbflXEvIk9P7xfgxvHh177bdeIVXCE7GNhxp1zOSG5ic+4Jzvg67bRSXD99ehURRoReBU
4MwLI+b7/y4iccnkJmkirxlbOIFZ+j6sbZE9D+ZrwNNbAUlMp3AfqzgoG6MqpGiX0MA8pFZFTmqZ
r6fZg41XGiFKCe3iPN4XuhopkX5LoEj7qsRORj9TmWksR499amA6n0NKCG0pPtNZlZRsmq8SnkOe
cwOZZANMZhHdQZ43M/LMu1gPDPWbkvWgEABg5jvIHzPf/245Kqsetwx9CRua2YFB5chFKnx8Gq/p
cESgudPNHnKu5GBCCTsgGnmzQm+5A6tTvY6F/E4k9pQFfpe8jykFEBM5A35ItJRX3tlo+HQKGdn6
woihxIAe+nCeGRsctBTYhHvc0qeLsaVL+F+Cama+bjp2gIyzF+tiiDyiKZZu+EZ1fIHWm8Xr6h6R
82S1/3PqSt3u5ir9cAWeONn3S16DQ2nszIRFPdquGqVZ8pN6Eel7ygFhBuMowim/CDByg3uknko5
zrgfCU4CbsVtpnxlQVuEmLZWIN0xwXFWdG31eysP6AuiBLDD4smgeM1XODnGGJOH9osEAHo3LAAV
2C4DFnj9rChdifZq+G366OF7yaS62dZtgc4BV6pl4MUYQD0DqIjROv4wXmF4ZIRtCuqCHGMNeb+V
CRfl/w5y8BZAEGhCNGBvK85jtk59SuFt7MOwJLfwqtIgL/xGvMM0IPdsLppXBtll14mLugSQzxRT
22tXk/cYxXzlmM6Erw0yKdNTRan+NsoJSt+UKkfBTeYvpDafA0XQCqM8cYc4TQKk6jqYAl0XeYo2
C7gSpPv6TOwWW1vZ5+bEdSQyhvj+wr5YJ0YHv9UdjCuVjyS8vTjEvy+nvvLxUwozEk2M91wkH29q
3rPv6XSRItZWDgYIEwHstL4i0KbY4gJ8PciTaUKSFiDb+OMXS93pdqO3wCib8FJHyao+rFQ9d4tY
6TjrEg57bgEww6er1b6lwpfHp1jWGrmO8N+9uoMPMe8NOkNccpnhCmCcsMrJjkPYmO8YCAcxyYC4
Rw6WDORV8xgLDb6DqYHDQDD8TLxbJv7SO8Gj3l7MqUbcT5wIGzAYm5vBrPYPvaduhrgGRZDueU+7
zUGnLMv8jDOQvGUMgm/6qL2qr7ycf16jrcYtCiNhpTgALbxGtJj0wVO2MUnSG42l4i1nCGSjnyqY
1b/iC7tlnMhKfr3BO9ZIwqyxIt8OW5P9Jm+W91esc6tIog3z0d5gZ89d5JZKz4JgDzu73TfBvZXs
PeLZQ/UUa0B2zGZu6Vos5QbdbsfC5jm0jlSCOr9J8m2g+gOyxhToQ78oCsJSLTfOzK+vxIiFXw6u
Gzbp/jPQ5iUaKjxfBr1R0QJH0E4nmXRadZKtjVw+MaGJBC6cSKF4MzYkGCTnYUROLU83ifmicXrY
PxLyeDBWB/mRUPE85PzpId2Y/q7D69j5NLdKoc8H7cO4wp2xa55kChdQNklsvxkZCbv+6P1OVCbg
DnEbzW5z1jQKhb1K6HA/O7gKT8p/z91dzf5ZGHHjRBAm/mv1r8F/JuJYU34ISH+rj6cH2TojsZRB
eu25QZ7r4wD5C0bi83twTyhat10LzmYGDFOSlXFsFvRw1dUa2xQ6rTwjhFiqCJGYpWlecow7ST8J
YUYbp7x5F4MYtyUyAK2qVS9ZkJY7q2MPj+qeOMB6WbWyEnDpc5SSDWX0T0KpxAKjo+Z0NEnubFKz
HnUyAbGenWBGLp/6ZxcmRvGhbH8ls5N5RZ54kTfmx0DCVEQp4jcQjo+X1tvn/JCYTIc9+KtDXSOk
53PD7QwDly0/5l7uWcQIldyPoH0BBflKkXmgriQ0tMlaXo4SAnyg7x25Glw8hTu/pq3GG4mUqNOX
Pt0M/mrVf5xOyyvfIE7JSjBgggBQMRHB2PWBWErf0bTC3WB79r2YfXcB5oMDGkoWsy0MnkAgrDc3
hG+ti8ISiqe6IjIpAnmxJDKHCGPWTd21GabRbPVHAeSkvTPZXRFymiZaycI/luzBepzEGw7VrmxY
T+Kq1hkUHaRJ7a0V5E5PcbdYRjsAj3ZjiI38UVGVWZHP8AyyimsDHoQppvPZM0iv031orlDIDVR9
P3z1BrSyUcflQDbINxV9xnmfPjGMaS2bQl2dbW0el/VPaN2sroOfmfe3IIuqjNaK+gEvEgFFtkzV
YvSt7hNmD1VSGwcL39CNnbm+G5d/QUdPQYTYDpjl8xc5SkUGXqjPTYBmwSAhZW1BpCuUDPB2l5gs
N4yuwET45ciknffOSLHlZf4u11nS4mzcOTVDBJlHpztTp4tvbNmz06SGliR4K1ic2NuKt+b4L1Ek
vjHPMdny8YFu4ToOlnerF46JFFQugykBUWQno9rFlHfSvuFm5SJlJpBuUv4zErToDb8EdAfKWuGq
YXy79cnHxMQBqYncAvScBeQvnutZC+XlVj1uXnOAQXgvtTQUc2wsY/wfBQv2bJZ4prKuYXKkxBUL
VqRqMgTbmKQepmcMk3Nco4bDyNKWZa+n4sIzGIWicuJzPW1wjctN7n6mAPLB89F6F2ugV0QTasCq
Zj1vCDmXTpdL5aOPk8p0sHRDnpJQ3aOt6lHFfJtqQLbl9X6A02yvE0IRebHcD3Y3oILzivnt6I2Q
lcDfcT6cBnZDE/i2qR4mvprYdCxwkzkqsJehZtk8Hhs5XgptOOdXLq8KPHWNawPsoc1KS5MJvqV1
ohmZrb/Rb5y9GodmZs6UJsO39THCANYxgthdfEWSqw4DUsu51sShcoPDcoAEH91HGTfiYrgFUDt5
Td6xawHQ12Pc7hw2UFujlGKQyiH2esjLoRATxiRAJKOMPNu4NHnscG+Jf7occhi4cwB/jR2ptkmN
9knULEf23bAb1wubVFD7YSehzu43gsfrvCJBpScoPyVEySg3gEm17Nb2WCAUW/4eZNYKtUN4AyUE
WjYxeXawAoLHZUmb/eyWzmSs1iwt+8eAHlGu1RTuFyphpiyvZKEfzXeJuI3OdHyMLFj/ndp8ijfC
TkC/w6r6Y6KXoIrU6w1q2JazWDqfxoZcOMm4DgRRo028eNav3H3zCcMuRTk12+c5pTCSZzfrPudg
8vCdsZ+/5tDUHIBLVe6OLYLdp+BAfNAEc1kzI2TPaLTgTyAfHoevQQMiUctR5cNp1Iloh5OP7b1h
BwJ51BqVCMJZNFbS6wXf74KD4jFDgemoLuzxq5ebCfWyg4Lme2KD/8XmJQk25t/o5x/S5ZRZAXMg
gLPai7k3mclRzI6bN8VpWBiscmcCuCgbMqWQn9RPVuQfQgH/Q3TdRfhMz57y3s8c0zLtN9Sz+iU1
kjiuFR4X8/3GtbXhaWNbmCCv7IIEqIuFod7ESdvcRMW//Hletbi7DrJIWFGWzt60rt2QuqXoZgLl
x6B/hsQ9GU45WX3jKdCPIgaV6zB4hn0Xd4Uo0UHnAgS7qUsiyD14I0xSXfei03vChEaMHBbBuxfM
iqa8fQXc3afHqDxnq4iB2OGu0gaK5lx0PmZbEoPK2n849Y1mpMvc3YS+GwAsZi5HbTF26ZuqOyjO
bC/wRSco26xi3s/7JFbhmOEcTy9dw0WLXtF5u1gxPSZjgrSYQXyMhxG+x4/EKT1QAfodv6eodkcZ
anGc2RsKzsM1n4tpD7iuN557wZYswKpbtFEnFT5VvnKtAfWF0EWE7AFm3koF6L1qHf5PYYxNH2v+
RX2FkiFdhQ0RDuxfNDNNi/3cLPLut7jPSpZhxSxqWU6fOygxQKTa0DBt+KbOFGFrwj7iFlEarAib
nIR34oLTRPgO/M1X+e9t/T0T7zbX1yWeRMH0JOxCrvHSUnSdsf5iCjAn82yDHWTNWSMP83oSTZV2
3+MjprbuB1PlMfPNVaoJJbRSZ4lmxF3gVpfmvu7Qn4BeWxuwhtVzf+nw46rGsqPrtG58xAwJEz2y
ap1AlpzUZpWW4BSHvxQ//iMrq1K5Q2xhJ9ocQCS1jDw8blSdWowCk52iVCKidOvK5NPzwM7Hzm+G
0wbMTGoyO0Oi2nGPBjp6LZ8QPdHp8HQT1528goY68nY1n4KmKXU4M7Jm+joR6MH3RsX5jED3+Jtp
gDyB2GCajjlSBRVRCd+hRrKeUvd+IFnyjgRLFnljdbDGOc1OD/Xsx9jSfRd23DLRj1hvlX7rO6wt
siBJ7zAhlpiArnbD1rVt/p01j/F/1Sg6a7WUlgII35uiRSBkZhe0Emlb6679tW5oLwFe7dWx693e
siHoMtJHAttFKDaJ1NUidA5+QJX/ZnnoPiVqWkxEpMtfzbqA+NGgI5zNwtruE7R2Kn4aOOKSYBIm
7tNkqlJMwO3BpIlQdIqY/lKH/WdP2EJHc1YlC57nSEg6dRcuEHGQ1NSjdIlSjKjPvcdTGQ/A3k5+
V84ZnkuS1FnwZGb1l2yaj9ClhifWeHiIJdzlyWGiLOKtjbV2H30seX1Zm04SqlsZUlQqhrwqwusI
Z60c2fAMWiVQn541qQejA/tINtYs126zAXy2afcVJP12zwEF6xeo5XP5QTEZMJRqx6290XAEOfXX
6zvzn97bw94vtHpET//8REnLH5voA97rQK6St050kgNICNSsnD1Ro1shSPKs6nw8t9ppu4REPGjl
4j+xqX2sPFCBlPHUCM7fupltXgav21dWMdUvO81NQU6FziSdFn3uSv5/O6FA2mpFSSuxgBtbrXhN
2GyFSLy8nP49oEUe43DjwX9RDRKOuzCPoxSig1lPmQ5NMPlRo+TVCx4/JCcJlnKVojCajDEpFC3z
vGyBp2MeRAnd63Fzkk66+SMhH9u2AeWLi9qB5blj5Yo++gMKr+K9BJg+mtejU5d0dI2KFdKGqQIQ
hK2eEJDZEvdJoNM5fxlWtT6HMFttJ8v6dSFyRXtIaaWNioQ/LMcqF1t348LfcDRHy5C9DmW8N30n
fkbDs1kSTsMrWTgiUR9qOoGzvZdldo/NWO95ClBr7wkyEmiRirAIDLyyh49R+V9u27g8zXO7/o06
MpyPtXd8ilMxO5+2bIGoFER5lKHZBVxyrxWDe7zngeHJwvPZhDnAQTD+pxlfRjm1zLtl2vfhFDYc
FD+CKTG3g2VXwTzFmYF8K/Z6gKSLEP2NGGIm5vScHuMgFDyagwx3rWDH8SPLFUohdsBV5Umkvsd/
WGhE3x4F2H0MI5vYGGbv48gt+zt+avRc4WSn3BMUiljd7MrTjhFZg3slIDrpJK7PDs/iYSON2E7d
Qa/vdPxtr2+0zlWPN68PnY8HQd++C33+eVa7OwV0PN8wUei2BCGePoVySww9ZR/lkpw15PUEUrTP
zdjxU6XXRJlia1ulsY+cTkl74VQd7ofD9r2f6OVs0iMvxij5Od0cRMjOmfPJRwyTmVQcL4ogwevN
gOJdp2KtNJISLrAjxR5Oec1Q5opPRXHwUlOKo7zyDIo5QZHqO9k9Efjix0GBzbLxMYjccAZmGcOd
hhjRUHdsYQZhqAVFCYP8yVJx7UyHJN8IOB9zSlBpUOD+9rP3nIa0ydzUwbaEooCuHvgxtAVxF3GB
pkzMUs3L6gERSInup8+7VUr7+BOOFflLonzhkuLK+SGIXohuptT00OfXVYLT8Z9EqdhYlSNEnPGm
kMbk1cWy+ZS4ujfMCp336qN8TDL43VdA6WlFLYihEwoQ+QZrJ7SUYJYAQ7ZL2WsFYy5ncb+TGo6m
OiHxb+UF+TXFgka469x+xvSP/Fd8t1vqbSamyFnNgrMICkEwVzQYDsF64vfqF5mtKJVDWz5BNMRz
zIORiw9If2106eTNCG8FFnSATYOVJ8vCmolfZDIGRcKw4Y1HCk6XAh+rZn0+tBkShJRtDarlriLT
+KIaDFKPe9qmL6b/RO87wad+6qGxMHN3zupknjLqwGhAD7rIWkymDINsxuF5TjS5S7vC8t0qeB74
kDZ1dc9MZjkRdd+60oINE3MuqBY2qmiWjqadbfaADyjXvV+KNNymZpqi20v+9bGM0tcukKI6W/n4
eOESwD4mUdZ5zzBkc4BwHuis4RiB7+DsKSuDYMJIjKYiJyjEy0U47f+p9EBpvfPrybD5L7+J7DjJ
zl+oA2hH01XZFJUN5MJrzQgzEbKTHz5CyDOrVJ2IeMViB+98mSfvVhmXOIKmkhMVsRMGVOeekPdy
jZYTXLHZUcpJlUGhfLe0I0XEosepdIOr4h+8N9JHPPgroJxbrJXMv9NB8sPiQ4H/BKv6p5GUn3oK
wzIS6KvI3W6u47HLaPpfb2JAS/i16r4uWoEB//nouQ5Z1IQNIIQVWnC+m5eEGEp3mw1khlSPovmJ
3s6WghbQh2RBBOkLlt2N7mx8mZ9X9e89Mj/crOC1bWzeiZAkLEaqeDkWukrchmEllY8M3P7CdxQH
VgwaGxI5KmAXmV8Gw4gMXgtXl0KAdUT/aIwxT9HIpJSMlfXitrOTpWG4y0E5TKHhjqEpUwjcxJ0A
hVGaGnoEsphJrG0mi87FOZledCGj0wUohA1cseIHR0uw72PzIRtSjN6nDoL4UPfm+aFou1YwwBok
fdwK2+GuJJtW4gD5Rgh/7SBFShngoMB5abNR0j5XisKCdfRGxwIqBOw7CAA4hwrNziiVzvgNXJej
v1oQIcQefYH0/UaFsr/kdr6YRwbpzMccUbL0AucI6+pdvK3HoYikdfo5am902DGlvrlpb3o7PvhR
Xp1ZcYxEbbmLbSxJoYg7LRDxxhA+aS2hiGHln8HseMQwamhDQLhfA5X31QznAxDZOEt9ZmeUxDKg
uF2P+eZQTjET5yMvWEZdnejCdPpIASNc1X31KfgGLMBnUP/faqOAxW50qrm6vR9BHVRbvNy+5IWx
pd3BpwAJNqaHyaoJvCbnvEH+yqZk8kEBAyamw/XzE+Eo3LmiYiVbGlZPXeFNombwXNrok0h7lDXh
n0JYGJXl48bDysiGsvmX72z8CV3Jrh+TKvtq+xUQShHE//YudrLo0yCvNVdyvI+0dGiBF+ROnfP4
ymb1S8KqCCEpQFDqujFahOXmIXQXGiVg+shT9N5HZD9RBJ5H+x3nzEmZpevHjtqoJ+zRCdAta6iN
8nwmMlXKuhdi/OQghhAPKOxakOWXdC8K0Zk9yuaj+eHmHyWzk/HtSbr6xkzSq6VXletKM60mzwtE
VYmr02GJ41O2BYuMrx1CsmNhGpXx7FBO+qcGDNkgDudWtXZ26MWs1j/5/BiQcjAYTRtQ0+q/UISd
ShODl06ebWCbPRre2GawlwPkRa6pl0jqrNw0DkkyntO6d61lbky27U8KLA60WyYU2StYQ416g01g
1SHryAyW0s3pkEaMzs1WTTLAEBKsJ0+qBU0LFjR1McY+iLGq8UF0XAq4T65z8WE7+QcbsAmEzSt8
EjVnAz2AILmLKEoI+Y6Iwdxgt5bRyKqptnryxQ/7jOkeANcAIHZ9wA2ZAWgtVgkeZlpXuCHcok1R
S8c3MNQGBfKgBugdk7UY5Zs1fDr1BqEEf8pBBLMfHlXZpUprbL8XKa5UExgGznp513NbDsX6Qsug
F3Dyx032IpLCngvbvkj4MjlLkIweupCpyGzydBOwK8gVB0nTuFA+nOiUx5l0jTpssj3PJtC5Pi2x
Ec3bm/l+6X9ckEH38A08Eu1KhL2Y9CP0VnhD3MBp2FFysTpyN+fSVH+40G5D1Qtt+XyGRSm0EWcG
sU72w1KeL8WXD5Z/iefcKDe8zy5N4ee043aHEtb8er98aLW5BrXbwYGBF3HggB8SbsznlK5BDlcM
qK9Y/7wWozi0qESWeRAN/reKepJki0zmIE864MIxnAiy3CD4lpRLh0d0LhOYWNiHsuVVLsWRX77p
/W+UVyibdtjQF63L0cZ932yDSYBwJZwTGtGyLKOmh8F2eMVrRK1Xi/VWtH7UlOwwwj19dYS5ojDo
Abs1JE1V01vxBqzq1W1w0CF2y1ADy9SZfqVctGhr3u/Z1y5VlR9MwBaymGBVpfXcskK1yCNH9vrt
8Wz6nuT5hIrPRXZF4twSjcEnPkOkirrXofkn2BU39No2AcUELZY/zxuNR9sMcHQVQF1gKJb69lLk
B7iOAZ+1gCNI2lCQZ1/6fewKO8YrOvdAw9+sT8IO64O7EZN5xPMWhT6lAPLjgPHmnaMW5Iw31aYC
oVTyhLI5nqlbPPIiIF+NLtLUFEzgGqkJYgOx9ViKk3sixsQL1FL+3qEPUZX8oeTZG+I2V1bf3PLJ
ypzopXZRxGCLZX6lcegAMVeQSYacAq4/f9uNYw5H2bDjDlhOFRj/p+dIvih4ckyoYU8aNo22jNwf
qluHbXmMkp/epX5ABm5NAVoHK/XsE73TUFOfPLbRqJeAC3qKg4ICiPKPLLElc/hqtpt1iwC06AVf
1NBbdIyyvQPlQPV8UN3lcKLvceGjpgV87a7OMTi7iXVRx8nwaa+ZmT8RDFO2DMSK9hDI8Or+1QB2
xk3C1+iSuzYjJC/+op0CJqSoJ9dKaigLEHj9rSzU8dEonwu/mhjeIAZSirpxFdhdnmgBvU9L1j7y
XQHjpzjGnmxSL6X1OBewhE6nznlaZ2OH81qjaspSOS4n4QzlzkOPk2plNgBo/U25hpc34W2APa8U
xXwgJwdWVV9b2FFiFRp6OaNkzElnhioMBktc9E2VTIxihZ6uoKrGeaAs2OQmGB0ZUxW3QD/VR77Z
DuCv9bKth2QUeWHZUYF+Kq0AYpIevJI54El/GJy2nJjDVFpTqTRXHtvBq+58BmpI07FkwA+jrAOt
qZNK2xCeFoYFaGB4FF3i9n3wmJLmRFLGqwi33ETrNDyxcZQy99ZkoTP9n6demLzsXCLXVUrksSsC
JiX+6sbTF2rH0Fw1xe5GMZE38yBq1hguLIlbZh3Y1q+Gc1yrL2zV8KqvWJLn4G92zFqMr8sl+nlw
eJD3WR1ugvgASI1rfVUagZpJdcZidj5VSP84x0f1WtUd3FTYGajxSvC5L6Czys9DULoP/YXPBU5w
O/3Hg20BArP7cDnF8TfPZWneBPU4KO5/LCnS783sI0lk00/lEHxSNmgtDZrZOr/MwTruQxI370da
ic9Y1UbJQaPF25IS2lQPXx5pFNCnCca8YnuiQhfHCBPq7y9nOFaUb9jtHaK3g9HjiWftlI5mZzD6
npAhBsUvmobE/OZYTe30A5uFpGO2O5B+ufaMUJ3RRk0w0b49rsdytZmZE7vcEYUXYpGv95hgZX6k
MyUTxOcwfV1VdLdJkFKgk0RrPs3agjS3+yqF/pcHFm2ZkutpfQXEuxth3ab51AJ1snaT+rHjqzFn
QHSiEpepVq8ad7qNNY5O4JQWJEt5SFBz2O7jLTTAvSCN8ns7Z4MzuIgJzqVIbGNZvIHugrtTEPBp
VNa13zV6CRE0Kyx2vAoeP4dWaG91vokyKBCgYTo7z8ssMcMJtuja+UA7g2POykewlRg+3hrYo9Mr
ACBXj9xsg2bS1TItyyWGPwt5i1SuMzTbPNyBt/peTVbrLbVtIpkjHYCcCypBWbG6Y+QLTKzvNHrl
eqiuUMxKQdWkBjHnmsaTElQfpwxjs5FXZIlKVO3Ia2jNQOC0M/iVL0Phe8l5n1fV6idh1wjWdfgy
lnQ59OEfhv7x1nXWICycW1NxAz3CGC9Hi2CS/tA0Lo+dZoT2uAA88gozYv49tBVSJTJVGY8kQeRL
wLIIKxqStu8m4YsgQH8Zrr+vcVvqa6HxhH8giruY0TBJLmr9wiSwhC2vQ2gI8CYIg89jjjzVoYFp
JiXUD9voKVPIri1w5pHW4AKJpYSgkRoJqbH/gxZw0iltyeGZNq89+YZ+iTzoPJU/UnRZP/eZ9v07
kaKdqsvL0OrGrvWzy34ZDRDm8Zaf+kBoLnL+hqTtkutQfBOdoG9FA8cdaSBigkTwXfBIuk5rREX4
xWtBooD/QSO+EDNaZ1rGMelOh3tpIXPcYT49CHMfeeEkoorAx+WHqG+G34d6+lYrmtruByQ6b8Jm
sOSD1eTATsKX0zReUdjwk1VUBTPhhL7ufwuFePxYZfkomg/7vIr0VtYe5YHc5XSF99z3MdqqvgZq
Gn2Li99dFQBbCDG0n5IVeaMxR4qVzfJXNWPcwPOHaSulbgriDkbW732Epg3zguUJbYnm1cl1eKOK
nvLUmkgBoWI0+OK/yw1ZkpFaEr1iFgywCN3v6hp8QtmbCxa4ycWJixLpkAxURjoZLwPEfjo/jcJb
uETnqf2SIj28Id80bLdcrVsnRvtW8eg0QIh/tAy+f6QAnypZENsWZD0+5Bk/xYWRPxPLY2PzMt3S
KTjafYYOfBveI0okKSTfVNHJtae5bbl6qX2THs2BeKanDqTVnHzjn5lSlC9N9bOggaj8hAgMs4RH
m64TK0BZk2a3/stn3FzxMHbb4c5KRM+POO3UPfT8LsKkkl/q2zJtum19jkPTOE3qvRu4fG/Nlboh
QpD7G3B2/tYgKEFfNnotJ49uN4FXfhfuvjHuFjp5HDBXdzdI6eyj4MGDIrteYQZoumG7AVJM4b/w
w9v7n4AMeGhXEGJ7yFqTeX1TAUO4SUEucFeGhiDuiG+w2VELhwsPUURQBh/47ZlkfGkeyWc5e6EN
gQLCZEJhpspghd+93LvmSb+o3rWtmueWP3OS7cDOsDQiSGZ8n+0eilX9u6U/ly8ovXbwTkGWsRYl
DF2jAlblZ4swpcrGisYj5DjAWPfuKlQ7zdTiJkaNB2ZlZTLJxX3ZIDHYYI6WFM1/9ULlSex7tzde
I5s6bJZz7K+PIVWcxUuD+yHEUgQTvayhwSexhXKLGCFco+vhlEwIZnBVeQzevqt0ezAHGWxzSPN7
upHkQzDJZkPLJKvGBaFKjflNsfk6QjH4/ftVhN5x31MQUKnTFMS8XO6jYV3I1e6NRkVK7JHSvszs
htJoB2/Tf8cL/cypp6RYH+b1mgbopHZbTu5BHzfm7yYdSshnATH3ykhnpN6iZdTftGhVBoup3lFd
XUPFi7NmpJIhFg6XsF/vpS5aPhBn7j2ZSqZlHT9IjtqKxTAy5SBENYSCwytfLD+Bq+RTzfDrhdSz
mN13KgM+DHKzMnU4uyt0/qeCrPYvY8FXB6HchYkDrppVZ7kb3gP1hQWtvhtPNTknymyPWutmvqfA
UolYowP8nNzDAMOfZ8yCySK2PZ1LCdhc2Wj2VxAV5N4X4Z1KUWyueo4iey0MkuJ78PUy9vTkWOzy
M7Yko1lJ4FWCDoEE5DO14/N+bhKmxr2FogHjd6VDaQd2bV5sWkH4/FJOe0tNrjTc/AJL+jf9sP3/
lrLoo0J4Laal3lkt+sU2EB2475wm/47NeOEsiDUyFQUxg96BgtEYi6z5AfQWuHhjzFuc1TuS6s6R
xlLsuUPn9dKFJllrr4y8z1mh5FgY4+7xj+bD+6iTg99j/R63944X3FwopJ81t4Uwkce5wqVCz2b7
bxkZyCMBfSpESq35Lg0gfsOSpcCier/EnIwNiSH7P0frmgCnG3kyUF6EEzxy2jNkZnMHkfMzANqY
zLVqdhCt0gLpBAQtpl7IBvpb1QN2t7YPk7aYAMYbI6Q0+8BoTc6a49ixNL1fUQXMCCayHRRsWs3k
TKxo6EdamDEmeVtGfZntRGe+06qabGhFZJ4yriViawcVJK4HvXgT/mK/MYRVkgXw4YnIdgBGRxJW
UniCpD2u9EW6zAll3irXGWGp+Ys8UWNqWnybTYW+24VuXSwzF+GguIzSpW0ruxVQPXxc6Ijm8gY0
6shUyW4RrlJFqm9bLXFmESvk1k/uDhoEGpvRqzzRXwXzgQ5snvgKIA+/0MehMV24DVMzbLccEFXn
mzZ/d3Zh9imK5A7Id5a0zVKD/VfrnsvWjnjKOuIm2Sj6IYABsGse8GdUPoO7pll7n/UguO/oS06/
Tw4k+H1U0auLnYfmhgq3eXU6KvTIlMU=
`pragma protect end_protected
