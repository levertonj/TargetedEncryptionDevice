// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
n0AaVWhNOHMyCY5k9xULNKubGfhCkWKHR+2X5UewiCZljVM0C5H1N+k4Eaq94jW7oR7x/TS4NWv2
u8i6uRjh0k38Nci3opB4oTXOGPblaNbtMehpJbG5jMd7XF5QJ/HNFFd5k7eR7DIkZVw10QdTziED
9JaqF7K2sxFST0RT8DMGvJxrAUBmEpNj5FLDSC1AQO2zIcfUEw25tkgebCyegn9k3sFEIdPkALmr
HEI/4pHcZvcm7OncOLbkOwbIGisVVa6fuOMXKjhj5gweuU0v1QUx6VsnrouFSx5E4pfAUQjlrdvC
8C7jdSljY/7tzI8UNgtU+xTBrXZ4LNff09IPmw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
DiZdHQVsD0AaZFGqGIG4YoberPEG/lg4eBT645ar943BWzqEB/zzugW1Z6QJMw8xOHotNlGRiPhY
QOb4L7FtaFKw//GJIHBibv0+vzIyUoNMMe1QICRoL7ashAgCBKRDZrA8JPz/gfyZwotDwgTGM1Wu
WRc/Q8AfT6wkXV3BdQlscp2R6bdYRvVaukuhMIJa8mLdPOIvCinrczM7boj9OHbdPocxCHlEbGbe
62/6gV9jhrJdnYhdKdD90a5MBY33uoQabf3eOzOSRhxgiIfwc0BO9M3absuP3vSfsPVAOSqevuUB
E/LfSbXB/Mxaj04YM3BO0iqpoIXqS9IMo1wWbfnIFWWCzAbsRIJ4F1xU/KuvlZp2L9ychD4szSzN
1/s+1aoFjc6Kfzqhj2QNgZKKtuUCSsN6b31P874P5znzeyejA5TPZ6jKPFoUU226wk2V8gyKQuuk
HrKbnp8q6IWwsWEtQKt5CNNuk9sC6Ep3QXaB/hPpub/PrH9LFOtkEfQi2cGqqBDthYDsk/mAs033
0zxj0ABaX4b6IUoGrdcnVewjba6VsKBkyH79IKWpzgm9WVgdolIKlCptDcZcb1CBbEPlo4eNm8lr
jEb7BsQ6wa8qv/5nyr5gOfUrYUrbtWaMso2NUa1nLEvm+W/qn4a4TYI81CRUK+y+YMW0jpSdyo6J
CRYbDyGZrPkNviTVFhoQFIz2jFdIa+pXnpi9F4uwWCYq7oeGtGgAgRzbnXusWMsIA3drFX9x3BJG
/2XZ01/FEJ4rJbhtE7A9hKKMFXrqguN9RXwWKlGwvF7acKM/+/g9PoFFN8q6+nm3T4zDtZjXLLfS
hl6bn+uuuRIWdcLaZ4WQwz2gL2aR8j6KuIdkWNIHiT932vOejPDn64zLOCbSlEgBtsLNzQ8r8Dg3
9jvze6FmnbZ5/8wkkUVdVnM11zZWhI5Qk9Yuuy7nIjtotlqNRoPptbOK2oxwzypjsZEYsKxUGrH3
NuQBKPig/ocW4Vy4gnu//IZaxfWPLZPcPwjzHoM4x9m6WNc3YmW6mhlXLqmn7r3+P6Ca0tFZ81DP
5g65YWTtFn9zZA6l6TALSqSU92wjANnYr1iQ5kOy9+Pk3I8pfMFFSO4W4mLppzfoEbXYvBvUKjB5
qtLWBLX8Ys7ktT9CZTPN5URQILmHIYzMBPsM8DSjA62f6LLpM+BZx3Kz1awQPhyEy/QMCzjTArHD
9EtZMgUK+PFnsk7W7gWEyAQ53rWA+lZ7MZ4uoXFNnpB4y5+znuQOciRdc7c+R4GaKi9NAHzFMFrp
qiwUWOLmMvEd39A1kU5lDFQ31Ntk7qVg4hDxCeDK6fSPSHt96yWnDlVi76mOLFQK+8/D+zf1yeXi
GTJ/rWJF0BhqAL4QFVx/X+sgWvcpw81B2iCjAQ1fLt1KGxp+bmQNVaw05Gf6aFpNmnbtcWMsWA2N
4AxDNB/bypJtfMxDL9f1DGlMUBo/wkupa+gyVPvtnmBYmDPMI+HI6gyOSb78QC8fOqLDLNA/bHvD
mSc1jgK+xhf3UD6NJryFrlIvsM56fAZUrDc1GigW8J+8Ak2mYsNSgNSuvEiedv7ZP5NZrujvm5Gw
0bI+D/6zFla8RT3DJLx0oO/peNBrGxPS3TUD/y+9bIBsI76TYzhgOr2mMUZO0KLM1U0qFQmeftEh
Jzykp87NtdcmPtJXV3ByQqmaG9P/y9x2O4aK5UjInINt/2R26XuJ5fR7G5tvHQyTNsTyFf6viaW+
+CA8KZM+fhe04YukIMBDP6TzjsEg8j7awdJswJoVme37/EPAHCC75pUR/bm+qbn8/Lx0J+XnUyW8
x12RUyszZ9estMH0NhHveocmdkyPZvXPV3tLQptQNr11f4avjcH1h8HRgcdj0H2AAj+MsyISdGV+
vPkg0+qwHl+ik0Dvg5XqUBDXQ8qnSZKIjj4NuQ+6RTDaPPNhiHafcqOybV5YqJjB30qeNBm00duI
+Wm2FeW/DUoCER0lVKSkgzp29PjdAOFmbQwU5AH3YX/P0UKeyliNc+6Lg/rnSt+CrBQVq8LCvWpw
4XDChmvO2rt9zr2iIgIOEvP9YRqsxNDmWSSPSUyv8/2+C4Yct+Xab5VEUrZbNDHDyDbbUCV+5h4x
zVlPTEGai+YBG5Ky/nbU6QVltT0L/GBs+Ce/EWjXJKexQgN7IYIR3yReTV8AIpnbetxNmgmVgXPG
I/Jb1n0AyILxfTqbkPP0URxRdLAWF5eLmP7QrQ7v26b5UfY7u0OySbiI17VU5zmoQu/0+YRSepdN
222PF8GypGmLzpyFNpsq2BVsmybBN7enuyxSGyHDhbliXHRcmmAHZGMI3HlkBK9ObjwxSwhx94U2
ChGXmhPQNa4qdCwArL7/DR7zEkjXv9Gw1SDgZdrrzaXM3wMt5YHFAshJVFRFPTZLLYQL18HF2cul
Zzk8ej68kqI0s+XP/rN3KtIw3CKYau5Hr5l2RXqQ98fnd26x8DYa5TFxheHBf3lq4VC7ZDrHaCdo
i3VBVC3CP8Qytcjds4fEtysLYuz4oZ7vyK3B76KygLa9aj0bwhKn6a47yIxj4SfaCeB/2Xl+9GNi
zvXl1fgZJp+s7Crm113k6NnsSq7RzWzETZ6jxd0kss3lDMkX4jn6ElCZh8WyFKsn8zXrS8S78dF+
atCWIFRMhZ+/EKGNTB/wgCTfwmohlR1mRsjqRwP++3DHmc4KaM6Go9rvtS0b4OGReXP5JaSdV3cH
zRNRp0qcE0h1QqY8D31jM3Qcn0Arzf3ectNR1oUZ3bihyyJSL1hkMdQAxd2bWR8YakEozeBYqDQZ
QqrGHw5mm1PKcpAJf4CVRBel33Qa1M1jfKzEXIfRLjMHkk4sEgxxAyslJLvIXgR0CXeIBl6N4KHF
Eoe86FCIVayDvddaWzvWNH8cbBoyfUTwF6u88VvW6/zdM8C3m0F0g4YkKf4LgdYlfPxbn03gE0kM
F0wKeOpptIXrkBv/Ti0iqHCpH5AyDrpi756cX/8FHpq2/hWp54eJcgjniKh2ejuDo5ApGKvsuRk/
6fX68ik2lsN9a9si7pHCf0D9RSX24bsAbrVDF1kbHBpMe0HxAt7TSDNhI9dJ1zSe0izGYwbvPrxt
/0Vl0QPGylAzB5dREL+ChJR9ySUVfCPY309VLSjSgiM6Z1IrP9IgwzeCbWxDKfvhmeKg9Ov9IItC
hX8YwJkqORZ2jjk/RG6nuRYtBwq7+OOog1HVyU1+uh5iCgFHwiJvaFnOuHRZ3ff6BkvAOue+7uYV
WnWG2a1N0zCZtZsb3ulNndZqJ0dnIeH8Epse6qA0/bOpgz5bGqDFhB4ytRsJ5QYwZcwV5OQpjnfi
UdUYs+OfE55iuzA2WkVm93D6xxd2FOlgaPN3SItUpyBgKsUaD1zFKOppTSBv3x6pqSPgS5c+8mXV
SAKMea952Wrjgl4VEJyW8b8E38QuazxolPc2dyPtHzLCp9FYgrcNs+6r7A22McVPwV8B1k2fVj72
/ucwBvkbGsr76tw4Ve1HxPi19bmCxybK5V0++sIo1Y9IcewQ/8Cd2YRj5JgDrtWZs1Je1f3WRMoS
Bvn+5SfDgNA7u0iB4jwKTJ7FDgK6sJtz08co/Ge1Jy2gNQSwswMc4iGij1DvwUJrh1ArvBaKFVLQ
m39HG5iVToOBnncXlKpgMo24cwN8T+RDfTyGqU3E8N1/uEJ3zSHYCgjq+m9ASqW7+zudjkz1Y0tO
47RIa+GVGRNBiLt233VdqkcIzevL3EM/RWEPZGEdPARPqM0/4TCsRq8XPGQBcqOJIAv17dxC1MaB
G+KZ5hpmNQFssDOEOoEgkc06v6rVfM3okvxC994t2Y0IRxbvc+IGHL2EkfbhGQ9nJg9P2vFsPyuA
gfJSbhiGjta9IV+xQhMfCVKRWytQ9zFaa5N2sNgYEF89a2EV2OQdP+MantYqJrzwG2jjZCU4I1pp
6UI8twi65IwRJid0JZhN9QwYe+HtHrJGKD9Mb6sFZT35sTRFP9Uff1tTz5v8FR/QOhAO1ziOiNZU
RcY8vAk3RpTzhn/xfsrYq+bwQOi6FxyoQlvRsnZBTDv6KyleYF8zGPnvfjE6zNJfOw7t+P4DmZkq
9ynJhRIJn0K4jHdQtOvPoV0nMkLts9jVYLQyWG06Zd13JE++6G0sQpqr3ClDq8Mw7gDvLbchF5mS
myWBW8TznneRoh2iannCrLv4YnegszuTreupVJCXwPLp5i6EuzqoU4mx9ccQhIrCF927A3e5qOwu
JeqAI7kJxj1d5HwQbXE6HC+wjyrPKlosgTV1PWd/KjN6p0jEgVw82LIz6Jxe0DA8Iaru4XqbqBwH
NRJ0waoAq8EWAt4CcqPyxnYZDoZCe+zIoPV4XmcNUtwQeQJ4HLV8qKl39uZI3C0708xjwRV7MTWF
vm64mGzwfTu9p2O3Qmx4LxkX6JVcmOo7EYx4AmjFiIJD6uJY8EdGcySjPv72yE6Fkv7c+vDa++Aj
qJSNfb2SeOzzXdsI3qxufptzk5pHv+565ueaHkVouknOmsDy2y93IIu/sKPGJcCRZ+mq+NYtot3Z
5xsf75ttp+7eT7TRDwTODWY7F1BvrECtBKjWyCt0DIkJVBBQ4w9Gs9n8b1CiwCEvq37FU05eUbNF
liNPM7p9RXP93ZKDivwVrvz88XaOVBGuqWALG/czW018ty3OUemwoSKTYxbFhHpgCkK7BFzZB1gQ
BPwtEAu6ju8pGhbmAV4k4VTQRrQiIEXm9BsEBFVk6pUHQR3WhiMo7eWR4AGDRLgF5PfDsZx+zALY
3RrSP8Ig7xcZGxaYUkBsvi5saLEWfKGlTZ1MUHPdnn+047Jcp9TeevJjeCA/frbPRC05f2vtjD/L
bctWuPw5gNxx7ld4EeP/5bFtQD1aBdxD/QgTG8znyQOYE9nXvupYPOBEyhOjjIVyY+IWZcaJB/rV
NAD3Bs7N1x0jKAul5KUk/t8DXIBrtHGxukoQH9hPPYAlOB7BELH/cCn8xIkM8As/1Lcb7h4EUyTG
MsAkeWOKTbjcat7tcwcOogAdIkxVm0ii1KrEuyJhDV46YwOxCka0SOj0vyt5+jnTp4PI5joRtHEE
M7/2wl5r/1KNZeHOJusAftACMCOMQPmWN20nYlS5NvL2ZKBZTkqPSwk5Imhud6eqGvRcGd1TcKnc
oGDVZIQupDUkC4IWrojfKHCwdZHavS7tq6W/67HJXXPX7Saq37nquGf6nf5FofkI/p6MN6RAxvls
RUIe/cifnBNtsY/9w50yf/JxL8VTS1pPmGoCyF8W8iK2xUN4Co+v/6L7x6XEUsCcSXySOIUgNOmW
OQ3SO4DOJ7UU4uVhTbPvw6sWyYN5I5wZ0BGLaBzUAx9YdDsg6HalFZ4tCqwiE1mPY4rHGKkwfXc7
x1zFMeufp9WktbSszECvZjdZqviQtvqPI23SzhLJ3kvIz08qsO6VoXxkYoEB54w/Z2vdkfnqUMKI
Z/7QtQw90raTXBhJqaer3eI2TzrCDDvMB4SG4emlVBy5FGILzWMaxTxgG6lJWRTDbcbBDEbF1mV1
mh28nXs18Ib1Pi/rGWQXi4EScvg7KjXaHNqMbN8myb4buj9GaZ1JE/n9+emJyk3nGXdtAmpGpl6U
qZuvNN05dDVnK2UuJyCOLLDhreHkxc2o66lOPSTbi3ojIxH6tV6YhUYWWjITgg9yhWHJwW+ig0U7
W0eKyxuIPH26TgMSzzbiM1+01anBT5xzTRs/Z8f0lE8NUMz0cW1CoKpQNFkaO0k/r8CgxNDhw/ck
96sCWSKGkmvZUECaYB2zufl1s5/aFdnpAuvHhnNfg3oTdLikEZPxdgsiKRSnaZjE7R1WQbSWHqq1
jrkj8ym5u7sqh0GVXGpJAVq1Rh5td+Do9I7HirqxKMzLz+QQv+eUwtpuZtOoYX6lNoO2jG3bDb0/
WEs7LV0qxGgfC5qJv+UEv0DmGiDsle3I2M3PZjwHKCCvGu4/jj69d1pki2DMurqrD8/75dXxdju0
HFwLYN6cYIkW+ZvkZ5vY9yIdodIuwg2n3kGqMhSC1XVJA3h0DHaySzuap2iBkLwTo6GBDk8dERtn
tE5jS3+i01xLPt59i6uERffK78L7NEOqDwMnektbN/Qx6En6USqC8+zUPhR586vdazyiJ3Hp5guT
cfyYd2aJwDGSf2ocHGIC/xjUTUyUnFbiKmLSMI1+yQ26wUh+QYVJlnZd+1XvG4Skt1bfs4N++Rm3
0eAsIRIVMyQLQhJuAjzmVGDYM+h8hlHSt1yWpCOora01ZFkSQSuDCFP2oxMGt8DsqajEN+yeTLj9
m76Q8A5DQUfFQKtKqyIHC5LEpyWYyYVI7fLHcNhQKEE+sUaH9yIlO2i8UMIDNIvk8RlR4jCFMiAv
F22BOlyBND7cAeLvDT7uuMWHUBCyKt4xWm1+U4WibcpRVxByahjU5nT5iBreUI4QurM50S87UQjR
52FlHoNDgYYEKdZoVDBAycp+apUso6TXYWNsvMvngRdaWXMK+6ITwOvs00mOIlawshKMzjLd5J87
QKHADXCT3EXjhmKCMuAJvh9ZJ7cp7xEbvJgOBiD98+WgzLWjwtqCn5R1sC2JgmTfFNa33Sims6yZ
KQ6IQKjcPl+Lr6nAUMy22G41FxuI4sLtzXFnz0S3gLNNMHpShGJgffoOvp5FcRnmg1Vrxgoscw8g
sq/makSpgBzgTO+f8za1rFr3/icyiyriP90TSavDjArYaoQZXkQW1IYwgF8s0LttL2u/IPGMl0uW
54yCQ/Lq1wYfWPZxP4fgGMnXOmjJym92OO7miBenLPtDfAyp5eek0716Ifz0v1aVge/yKTyvwhXs
2dvW60y7uC0OgLw/DyC8v0fhUBu8ag00Qy6ZEjLdqFuUahLx3+8jx7279TNWPuMrstCCU12jiJdl
kzk7Kn/w461rG0ca8/bMuOTYICtaP8m4Xh62xop8ybLI1mo2vh0THiHuAFRU1sGpS+HSZ1pYsOb7
6MUWKIaIpvsooS36n1hiPB4/J+Z0PNy8ypKBt+IyWZRfPP2eKNP9piKo8PA+OXTj17IWdhFiFm8a
Ahs5r4wnKDL2QjuSV/V3M3sBNV2P9N3/0Oj3Nieem5AYeY9pLhpmDgWl5zPT8Rdc72G6bHRYWHrM
0WPTXxcJ7upL/o7hvcqOxsVRAiArb6u5QPaNR80BzlmTYfJf/yZoh2PalTSCBS7Ck3tLzekqKddj
4MpKR4iEXmgmlkmyIjv1zW9QrIKEU2wpcXeS3ZuWTS5ZSIGt0cS1F6FoQBekjVxGSADNyF1MtVUj
W51H3ip3hDg8xRxveoMCRIWCa76uGHCix471bw3D5+Z4FGWfZMmbexpNHQNk8xYxXzEUBOCiR/xP
+Huwk7GHLu/gppRj5VOh0LiziYLmHsYPalCdihRsWb+yhYml81MEBte6nrucXEqc61dJcBVPhxQ1
tpUR6OR8D2vmZIf+siQNPWaNta1SKjeqXAeF1tNmN0lbtZMHgNFWV+xg23u2jxCGv8AGF+vSMfB4
0l33D4RFUlNy7NtRJcpHFzM1bdl2BbFOHIyDoqfU3CgNfIcMf/guN1U8j/cm363+H2poahQ4zgNS
UAJhnJznjrBlBO7nj0jI42d466q66K3jB7cH6NJTd6mjbYG7Y5KgoiPg9im0msghcVd8TOrfKkBh
qlxz+MUkbAVhEGoDitQzZXTAAxbCmjAO1ZEl+cQLchf/w0abbadscVZQNI16To/cK2qsEiunCHnc
X3YX1EXdfqajZqHSn4oq72OoDE0enP5YikJ9DK/seB8Tdss4GHFVKGI0nAsdltFy9l6ekPSWrv8F
EkudjTjT6v4Jl9LsAU0jak0w1tZ82pgrjxlQqQ/THg0t2i8UB0gYSfpnbXRlKuy0dXpQI7DUk4Az
xuAQq06glQx1aSSyWb5VVZezh4Kr+YlPxeHzrEIgeM3ESo6sDKyp0j6gHv0BkoLouPVBCobc1I8P
76q4P7gpbreVHTEc/HkNepJhsjeFNli1z3HWrWpa9gAy2yByIyGQnVtJwmSMVcRD3zHVld8FK4sX
AsDu6+frDtGeEeGRzmxfuQZLzn49DRR3HzJ1PuRynoXCEYydEYtNzsNRPTg7kw1WvoXBYSOK4YvB
TwvYvtY8ZJ3khPj1h5iF/LI6FdErdEmwYmRgAp7G06K4C44OYZY34bOnD0+mrJyeqzc1q32MAiSw
DLpdbibz192fFInpc7X54j2LX1xkJsOtja9ALeEAxYPQPIS7af4iWGahofGTsQSrnc0dYSgGrnyf
9DV3lD/sGQ47SaVi+THCmuQbwChppVtN/ntTNWvH/VGbtWjotz2cVR9xjGIlou1+O+NA0mCbVJMQ
Q5Xe/uIWjSAhkAJa60lHePhflBLAnnnSeDd6wcyUYQzpu3d7l2tyCgC9josjhecm9pMWOmkofQCQ
Hr5Zna2GKyoR+DscwDyGMqN7/C/F1uaXJyFqdsArqIB8FQycVKZcUtd20enNFFXBpz68lp75YIwD
mW+zuJ22AKl1qeLiw9/1wLgRUiZdkSHLK1Ti3RbtZeuV1ziX5MhiZLyCo6WMtX2hbppojQbCMdEp
IY7o9mSzzAKdf+QEqwTO51JbUClTYDC6fSQ+pIwhcWAxhGuSaf0SOKDvSKuCLnFWdtrHw+/BMDK0
+PmRB0as6xx6tMk1svSNvi2lYrMflWO0th/StbPcxSnCLgXO1wDnv2tsIxT0e38aHBL/1OGhfc35
0tLEwlHwG1TbxIr+sZp1PzMBWf1kAbvVFcvnAqIgLPRR4nQB/7ci8PsHl8bnOf8C79A4rN8J/IuA
oFGAPvkOOkKfxHH/LK3beMq8p+npwyYXmMshmDXNOHDCwuiUbLhH1Fp2XcJJCxEb+8JOel27TUqj
JiFcRD1UAeur1/RsPy6LLcErYiXITF7PiPDH29vBKuzt/NdngLnwpQePuoB3E4Icwv4lYqj/wiVt
akWArvvPWNFnnjX0R7q9bW7LwYV2jRXup5h8MV5lxYFKQBSK45Y9N841bVV/EnvIHISn7MRQN7Hq
mkumDTphuO+GSrQlEUfn/VYON0EHKeleUhGOWa2vqX5veYCPWRNw3Wpa/tUZQuX2rPsHkG5wvdfq
2IN+x83ILgBDfMXbvh1c968HycCEN9zkTNAxCRMbYdHNrSOxc0ow236jQyJNsYRtyOwpYFQDw4k8
SHCNyTwMyuNvFPkxcmGdjlyU065bM3rNAB1fejRzbOKJLYuuuAsKEpRc5VVtPaqubZfp+NB0fl9s
UKQLRbs7xmAUsJtFAY0MgyaRrJkgA+fEFFZjIEnNLxrNkG9y29TyEcakd1CVQ062j8SYQgzMKyfq
9zdV0g6FSganhSGN9DBjEQtj5vgozkvsYGmTCUGURYJ6/OExx86fZ+5wIYd2eERyjPTpF3XW4cxM
msUoeSZrjyE8yzV7RT0D5QUYEofU1SVWPwKOCn0Xgt81VJyLOckoaYqMnNUCbLnPe2bx54LjD1tk
OGHPEGxSoPXcIZI8luvgoSOyPQQ2CzWFzg86y1AEpyjukald6N2Yd7L1rUvhrY6tE5ZHiBrE7hz7
oCWbfgj4P4aW2iUKbeuHzMoXMKyKw6eW92Ta7Pq98ddIzwbqwpFMAf7/QraSFzoxuzuR/Qqy7Lym
sWTi9OkYPV4RKrsUMzVo4As6WPBmRf13Syho0Dqp0lC+tY5SwrjZFSoZ++SxWUQOm3XRNTcRG87c
dPTWAQLJnQEivWJkjmhkxdpk2Z8ibo8bq7b5P13QHFCRDLboW8MAWCEBKfQ5z/NisABSSv8hBWti
ufr6vY4XIrxrNMt0xjd8VPkI8lnV34P0sobstlbEtjmf61G4apXl8l22G2cRXRPpmQpNI5zYxhHm
C/E8NdKXl7DqO+qmZL/+S2n+lLv0wjuBIGCYDuwCwXtcTdmHnI6hBxvERaT0XhsSgDtr8f8dC6t8
Iwai/Dj8/fuDYeNhPBgL84vh5BZwkSfuIrtlZ9Uc6CgOJL0vlrqnzS1AqB8yigJKGS4Cwix8SCEz
4E4fzcwP24WhRy2De9AR4ulKNfetIJt23T63yQ+i9HaTM/3Zu53G7jF31pXQBp6VswSu4oBHZNDe
/PBumYQyyOQQC+7lVZPuqd5Gn4Tm6uB6iuwrruXyTg1/g3ir0topQmXMIrw4rfX6YCy0SFb2enzD
KPgCz7uQVIpYNg5AqZKGVDkMQEh4QRksqEqz4bG1oRzhhdl9wooelJP3/ZmKQP4Kd9JPNVoOEGGK
svX5/EyJx8XT5ZiYhZqMfZMtoHMkuCmKSLE4f6xRz9jQKmhPVcP8Mk3BfU7uplenUF+nun+EkzIS
nuHnnLCPLmTWVlmaHABQk80HwTdeThOqm7Selsg2s4hJyUb6iz5sDNhAcrce+ybouf6WsF2trUEY
i3Qp+Q08MxHAXzs1Rx47vlqUnuumKVrQXkCXBcfl6v2qD5HMtJ95D6H5BTpDaEPj7yLJhA/GVpR0
hTMgIXlG+I+/FudKlwZjpHWcRuWrp8snhhNKC365f69qUVm5JGEF/jaaSlMSo0saGtqfjKC1ZNXj
/TBCJ1WoOOsNRUZ47i/rOcKsvcZlVx0qMM9kAU6nm4JVszL/g0c6Cgpry7dU6XiIFmtpA4t2xl2u
y48+RzlF4sk+IZwx8aQgCLQNapN5vsDi62XwjQPUxO85u4Gw2waYNwltX8lylu4eLwwNERFOVFDV
C/IWUfqTO54TiIrW3dAAffYNEuMTK6W7bQUoOLklB//y/NG4iZdixbXC/bujco52AN4l7zr9XQI9
7p5jOwhmP8xBGayhyUQU7xMXAyuZXr66y3kYItU9Tn9UVg7poGMmAWU/CghNSXgsxWxG7RMbFVmV
oRsM72NK617Mz5jTdpx+9Xr1sa1fvcYcvM0x4E587vZZIquznz+xjc6vsgyMbs76ZR3ZZlbdRkPH
l+/JfL+Tc67MVuvDb05MaSmSuvXUM6dgxCGxhrAdehMYZviCt3lFe7Z6apoNJL5MkZ/ilx4kG7Cy
TxFztg4T+TbLwJFXFtjK4llrAwHlGAjuMnpE4DeDmgw7/761sNDbp9vk2qlhBev3ZeX40RxiaCh+
7zXRG5vP4N3OAFgSEQbOGGxiR/Gh0xcfqFQSXMXeFDquNDDt4XVMJu+/H9SSnm7J/hXYf0ENXWbc
zo25CsmAFAktAkIymdjSfEM37htX/xvt53k8SH4juhjfnpj4+ieIqPk1ckIj6TiYdNSKR6Rm35MD
Jc+nKLnsQ3SFrAH3joq3+fwcqRqppWpt+hpZHpSfzs/KmYKi55w8BJVrT8q1ULSvHc3axlJ/jKbE
vtr976cy/0AMAis/rOjr1uZOx2CFQiRuxUo6jjP2vpo0H46cFaBwdNf8yzoEPVLLNcZZbzVfOx5K
RZhOlrbtZhjRFYnLEIBsoycO8Yxzst4sn/8GQYhn7fUzz2gqeZgcfbivyGuqII8KQg72drqcBNeY
ttb62WX8a5hbwYzy4sKxwcgG3DMMLtSq31k2A+QiFFgROwZ/DBV71yh2rZsA77EaXdhUiOYdzqw2
hm3cPY6cowoXIpRvbSeK99pyV6yl+U/IYAh3KRV8rZAS3ir+atbWTQzMDf6eBNt/AROJE0p3qK7J
F7fsVXJ4jbi/SUcq3yBcQ4/NkLYySUWdxbHY46D6fW5o6LK+SUcAnX32QdNFrxun8OGdt1rqkQ8S
OA1mnLr7MPFancqIcoaji9y2JDCn0mbHBoXzwRy9Xkq37tiT3TxsvsbOpgBCbBl/pEAToSvJCvMC
EljxEQ8j2uG2U2gnDIBlm0+vI5yfOWyGznFzlij45L5/HnwyQu9Wes8i9/iFZFrGsjHWXbJdGU4L
mxSBJkUOHonEOMZCa93s39ISJDXgAOXqp05Lwx9md40wjbqwPAqg6AfSB/E50TzAUdIx2MlTjZ2c
P+IDtESTG5OhsPmbXjd7ixF0FObq5I+LRhyEYXEY50flhWIKC53S/IEm222Ulebtdmv0Wq04alN8
Z8SkdSd181l+wm/mpULZAXcs9TRLVMHrExeiHvmeite6SbdPzlT+6Tp2TPddVThf9ya5EqZlj68r
OXYTOFjzDHvvOQ8jPU57py/MO+NYVrbDcMxmrRTG6r+R8KvaUZ4gbkH7b2lrozyg9Mga3+bldgo5
Daabwp5slKXuKQK8dmIgbtXKB3t2gjZg59nXdO3tDH/88gU6FeeljfGjszp62/vxk0H9nBDyMfvC
S11r9G2V3VEUbZyCfM5dVkMc1Ynqydc/BqLSU5o9Bl5vEaKvLooBZG1+fdEt7bw6yrTrvIO0VvkB
unY6+LeNogYkdf8dSEPHoRu/2zsztKONmVwp/eYRmc8KP0MJAGZIT9NqGaAESlq+Rn6kA4fjjhxh
ESLm3hYLTffZ5jkwjq9xuAL46GAUOggqNDXC3vIy52WuxFzaXaEScyC2Muzex1xOJDk+Kj1Qvi2q
u0rEAvUKWPIDAmrTOt6FKF9uS9yMuga46TkMqpEZ/1VmYIBvUZh/aiDVh7k7lIwKTm/3TIxvLkDH
ilagmwgTUuVIefZI2pJsx0LFm74GZmIdju82hwaNfdQtHCtlXMjCD4k3WkLma2Nnx0p0/2h+Ckel
c11dxpYV3wHjAck9Ih2zqLDRyQegZd0+iXl2tqqYJ5E+eEMP/J6WQf0aGq/ZqvjRpNv2Wg5oL1bz
cuvIg6Q3wB0jA8vvyFpBzDxZ9+oMgBgrURMst/21BRSflnUXSt0s08YqzYM1FeO/qnPT0bBeFRiw
ZOYKBtm0UqBh0FQsrr+6RYwzLyH7RgwtuMKHvrovgVLwKM2JlNRw0kigkh9OW9phP+JEgVv5GlWI
uP+RMC0GM9pQLTrWbyyvzNUkHiwFfy4DrM1+rYtjXCHf9AaVVJLG0iOQswMtxa9oo42BfJB/SfZZ
1Pvj9GEpG3jFN88wpdXec7DI94IGNtAFCqp/pyP8+1xru8gF57hxXibgL/0cLi47/IHlxx4U8mAl
DgU2vSLuCF+NNZr1sozhfYw9lPImkD1t6+o1aWhihu61PYBjLRkDWHC3Pmj4gfawevhfSL1dQXOk
czNbuaLio3JnQAIxoq/URkZr++jszGdKfN9skNYz2YaEOp5fdKbcUK5PH4yzBb+v8u/Y/GPQUV5+
GC4xOX5oW1RDELpjFYnXkFRgsl3AMsGSv1xgP7GdVrqLGkEq8Rvhg1LXvQRdH7fYWptKmdEfqhte
bECt6X3ZItthe8DaoqW46QKS8uyUejK62EuJq0FB5xtRL5MV7RdGIco6rE3hOcY6N2EkGd2Napti
ooZJkJfGfGixVItdxK8guG7ErcIQ7l3NDkf5OFsSNAfHxkx4QK6a9SF7Yog5mAecMbbiSyBQIHKR
H+xwg5gwDIWAGHR2BRBwhLzRtqMT81FlKVuiyIG3dXIC9nxVnBwjJN/pGOlhctpBMKInX7t4KWrX
E2EUhZa0sLY/epwhURatzwi/36lEtzSLl/MR9HFuYdnM2go4mZmbZPm8bhzpE3/GhyfwP8MIO6hv
HFmYd58EiYsPOPZ6hPCc+ykLOYfikzNnkFb5uw/5n88/+rmicp8vTE/wLVhtLSSuNBWu0Rg5rpXa
EKpiVsFlbdx+rEVFHL9YqKpRH31K0Tpmy14yxD6vyb+ShlBQFsMFczYiRhWw5oSRrkGdtx7MCWdU
rT3LRvFyr3ZqLnfAz4MAVfnMKiO4BsotxuWULPHM0FktmPuyopP7/L6Z/tN3TMIPOUd9t3t89of8
RBEZTG6ZLK1gmvoRN647EPkW4McHOFocZuELD6/ZsLz8T5UgS66XGuAmLH/F9qz9bHTm/UldZqci
s5wFqv0o9UzSyrUA5m8hv8ZjGhXbckYNCKNEAw3dpPKjbHcBB+17eQ+BNyvK0aHPiCqD0jCSS2AC
iLFCKpydGr5J9YSS0KScL5bUEeU0+TmSvn7yzfT26z9whPQMbLa+tMLlM34gwbv0byG0/BQaVPzH
Xla5MGfoextDsP0SmbPSaOumspssakH8TZGWMA1Cs+h2f0gttt9gogtHUxZefkzt+bXwk/6O4d0J
98MFzQlCbRGb6zSLzxoGuE93deguIdx8mp1A5C/1WalaVH2ZDvw6dP5CR8zKZpgO//u3tSCIMsKf
+U/4VStAz2SXp/EP+ncMPAGS1Rjo0hwUXLMpXpRhsHAsqUSgb8tnX3yT70yRG1s2RdzzWzV2gxBC
bxXfHfYK2FKWfaDkGHXoHMkO0weGCjTJP8v9f4YMpjYM6pOpc9p/kCIE8+M9JmHk6YDaNwQa9+dI
6qd6jaexCl21+3D1t73q3CTlzQlbIi4OMoDRQTo8I9vQ4A5gcgJ9laalwBdIuRPJuwe0G2+iDiQb
pL9WuVQS+KGFzvzEHIj1pRspcd4Yu2x7SLn157GAjPLxEuL17Yow0kQi4cIpV5/w7In5lbw9SqPs
c3R1ln3ysmwgdPibuPgLJKXYdsSd9hWkFG8I+ZVfugCYTN2gwCi0RrPOCpcbp/4Uxdc5THOT16lT
/gQEd35Fm+Bbkd01Bamht00oD5wuCHOEBNMZVvMGtJAkVg8QTWravNJp+OYRCUpgklxhgFhYIM4y
uazBJCj4n/fi+JOb6UcKklFG18dxKPsPgKZ6EaV29b76EPbJcwYPEYnh6mw/QtDoxjZebj1qcBzu
8ZvdascIsS+f2uKvtehahpMc5epiHd20fdGfouDkocMAB+cu5Ecw39c70IVwRmWQlGQ3v134pkMU
qDxl0FrvtQXfUvrcWlVRiccdIfoznZWft4rL/xrvPt/7AwZ6Ifi8j+BZl+FFQbRfm25kZAOhSe8s
kxQIERv83mXce1hB3mI8dRud++5ApYL+YUi9ZDbnMOB8HB+AddgPAeOYFV/ZGYuoigL2bAV+/K4o
bbqreS9pweCb+YT1CV2W9N+tcVQtzZluBhZzzmYAvzaMQgp+ywzS/9Quh1RRemQFa9Dx48UQWqN/
xwU5eFq4cmKpEe0TLVx8RHvEZyBJaJHhQUgHHFoPkR1FXERXfbuPuRsbubUdR2wp3vfES2B2HYqu
JtlvIz7nO1tT8SWX5Ua00LSQb8o4l6tjpl8zVtOygJVYobphhJ4iDsfnsitGEO2UY9W23gtVeCLd
7yjptn/rWLoCKAwxgCCnTVHF4esv/7tBShB9wuFAByG+D/KXu23Y8i8c8pfHFU/oGEkb2Xe5HD9T
zNxF8H5GEJN52oGNGoPYmcuAW0RXD6xsvBak3EdUHmG8qeQ2AwUfarmbcmzdmJ936jcxHDIsMgnm
apw9q5/jRJHRBrSZ1bB80pI2ckG/MbxzLHsAU3BWIhz/ffnfYOqNLZ24rUN7tebQoNvugVvLotPc
N6Ybi+OkZrjOmJ4WF2mU/6DP3kTm7/w0RMtX1AxGvjKfAjOry6MFiZVd85ZuobEcwz4pmqgsN7SB
Ed3z9RNTqmBS2QcTcrKdJSw+QAlDFMnRplgEpDtYlH/jlVzq+tz+QH56AknpirPZzNCj16Za0bXg
j24MV9kmv8r/9zbWk0TifgQQZ83tT2km5HQ2/m4VmBFj+dJ/w1Sw9i8Hx+YPXWrhCeLObOxv85uW
AJ2xXppV4XblKgOssCG7nsd2v+PunrX6hoLcbSAs7w6ZFV2JXqNGTgANeSCldk6km0AoI23Hj0Wh
/KIc6g+qho17uP5KI0+owT0+h7iMUkkY3NNHw5o0q0uEM2e0z8g2quOKsb/l8rB6kjI1MVFFFOOs
jIObGbd5T6tEKqocTU04Utu4SaExS4Pb6FDmFMP3ghljDhgCEOPl8eo1CQqcsYThT5jX26ouJcmX
9d74o5SdcjVOvRFwvtwjeMV/p26cifKtVp/Bogch35yQ6qVRMFXkt5CvFtC7vNbnVIHrsZZcVHXT
RNact4E6jv4SPuFjw1B7C32akksHYRWVjlVDJNDOHNbFexcS1SapvEbUEimyEhzfM7wuM0i8hSqB
lNs4ZmP5i5ddMbeSWRdMNv/dT3k9N0LxJl70/onfII5f+sxSbVbEAm9YbjKn0mC5yeAPbnxJzDyK
as4VnUsfsQRH+892vKWyWKfGUFvKcUF7MRBtMhC8FebJt8pk9Dbdd91+5bexwm5JOR2EhpSs9Mq6
4QLcwk/1GSm7sujlx2/NdxL7Escpn5FUazNchQYDISYH6nk909TIjh+4a6fwpxcMLhDerEsssrR3
IYn+rsOWcXG8cDs/nGpceCwwOGUb5mwCB3XOP+yTNGWwnD3dWFA/yn1tgyBiQu1d8A/Xm26lg5sd
wobiiN+caYJyDAd/w9FbZjIzOR9Py5mDCWAAIUOa8HvP+tJKdDcJ8k1AWoTkeqc8uyrYxNQkRNx3
3l3xS3zX08yAOURTkFWRUdvRZy2T2p6fJWNQSlO6UiCPziXQ785nXVHvgfJWtYRRnZ6hdN4LbcF5
FPuGB77leTiUfJ5kH15+Az6GuIrb1kMzC8PNgAklJ++9326BderfaSyJLXqom1h7fRwCKixRTAj9
JTkZryYLOrdMoZccpkUDpcbu78O3+Pj3j6K8swp7nWC6GBeuO7A0D0hD/HlVeGfaWy0F+ocuhU2w
8gkG11eOqnvEzs3j+tOJ3UseRYlBi+VCZt34JZs4soKT1TIhmokFXKEYiyFhQ5gf9UKGkwkJpL0w
rD5+ip9KrZquD0rJwJNgrY1cmg7M8h1K2PhwFAr00l+B8jWxxchF+KNqc/Jb80GsuKCpDwwFXOaG
746elGd4At3BbUJ14bqPVFvCOZukEISIf/TdCyUpuHHw09B0uFYf0QllokxBpNWRBXSqAydT0aNL
4hGwRAeFpQR1mzpFFMNNEZ/gmTBaEgWlpraDXs/V6Xc4nnRZ1wSYHlrOPYlg+7XCz0r10nOaKY/V
Lr6khhweyz/qV3EkwALw7yLTf/9pKR40y+UYcMqkl5HY6MHxqUvpiKu4GvxsmFIV8b0n+XGLAArb
BVIf28o0ZuH4n0+Z+cxMnqZ4NR7POR+Ykd4MW2pOdKC8+2xlZbJmhPeTu3gWA0Ck6HZ89G5e9uED
R8dlYdW14q1hkCFCtdv1ecljGZb1FYAe+zBiE3hsXNzCzi4Nj1dZxa/zf9gQlkKOcUqlx3mDNtbs
0KXpFsvBnQha0OWmCkXMKZYlYWerJisNT0QfqGdQAty+5SrpwA3onFcWTIURy5meiah331LSY/VC
/fF1nNNSv021tm6gYml5WZaqcE8t1a2M5O+obB1V/CPBBRNyg6wkZymr8Y3KBG2iM1frtKQkRXDm
UnySuf8JnaGe+AjKVDwdcP2sYkEROMhvclDOC8zu+POsIV2ZwdRbv8wFdz/zfaV0rX3Pv90XsMmA
ceAOZB62zUO7oImBlJA1K8fG3uyRAF9uxss7glkPTFS+vMNZEOq7xvpheRwBVHSbEpF33Nd5XDJe
xq1yTvhrsqCGnhX+e9wJolFTv4XtB+ptcHozymNZdbu/Ae6H9pZnmAjwg68Sn6eTcb/fSutn4lBY
T4PWm3xPyPj1o/37PIuxYWvD1tmfA2uK+wWLUKYf1YpTzDICHtZrLOn/CIHFEhzscKQGAePXfRk1
3vIOs2OVjMfPK0LgZ/4nqbzmL7AjmAdf+d8DaHlhDempuewa3b2GiSw6BqGgRCmNAkO3tckM7tSE
GoKq5YQE3Gr5OHB39Qsmv9WJlzzhWph3IfaLSstwDu7L4qQl5Y/bgvnleHoMRE8jTpADwP11+HPS
L02BEf+SWyhdtkO3/QV79ggiPY93LKvwEPL1/XmPZQcqvvElMAtUJ8w0/o2S/d8G+tAoIgZesxkU
GYa2emGn03gDnmSlHMU2xRO++Rt3y/U3/9kjby50nRGCZdhXT0wg2l2Q6naSAe3FkevZSHzK31JF
0AOgxreIwl818SnSFJ8tJuzIiQWCai7xd3TqabWChi4SLR0PIA3hzvr8htlYTJ/6EMUJ6aE/DJyw
inONEc5q7AVdA62omwOCF0DSyDR2bikAH9FDvmsNRGDgSvQ73v47rp5cbcBuhQZI/Wzj0mksJe4n
tu3rqZPVI3Lg6ZYBC0a3z5Dv9qJy92hDr6UnTxshlK6sMtEW7cJNzrCaKeUS3Osf9SpcNo+EItE+
xDcYhZIXf2Mbj/Sg8dNmgE3ZumN9duMHKi5qhka55hlK+CBK5FZa0o0rQs89wCKRmB9N/MfiBC+O
R/kA6BthGc4P6qCk8jbTjovXgtIfkqoTVZ5B4BfrQvncbse5dRRlxwnwbOXouKxmLhbUCjHpugCx
T0v0vn0sH9VZvDt6awKAUe+Cb+WPuNf/tR2mIV2j4jTL1lwT6sHeqfAzXUhyLaVhvMEGs9UlTnnI
6L60m8JwN1zOmw62dGNB2cJJi/1y9MNThffGann8SIc8drMNlNYBL2MEeYjm0qwJu9BrP9vwKRs7
DuTBjEENupR0oTYQUPgli/Z6z49rVJN9X/WUAFfGHfk3HUxeo6tMX/dZoRqHcI+LB3Yhn7V+rL6q
iBIciVKUNFkAdtePqnDzusNSbbyUD4eZuw5hwHoT3kqgH2ORtYcT6znJjMCxylrx4+Xpb96Cp5li
X+umf9+bKbflA6Zf9sCPMGrHyQf5ssSEzMiJmkyN09LT4JwWrSqbRtoS4kTDfdgvUZiwiVuN3xaN
qfZM4erWbFMDyrBXE2rAPJivJTgkgcMS8W5k0bK8/btJm7ZIJ/cGHw/4BWRy5EZPI04n0CVy1Kam
9rrTgEmc8m9LHTlax7odjbCnoUQ/Ix91MEFKpF5SvFdtIl7NQorcaJUXYKi5gDm0Vq34uWhp/Hds
5Cj+wFH7qWdH+q3Gwtr0IbxKVOBEjGW9xAlMushfwofBOSWK84wKft5kSi+ZLk9Bgn+aGU6bHMtR
5aLt/RIdecQDWomlEvsz+yqyAREIAavNYcbeCY9GG9fCqJhI4SDQdGo58669xJEPGW47OYCWQuD1
WyjxgSiLy0gV6ibX1NuJZ+VcWBpkAWg2PtN1mRtCSjU2dxuutbNye4KHlcOZT3d0lIpnbpE+m++W
HcNduTpKOLIuXXRuA8kMye46X/p2EfJ20Zn1ZzxuYTD3GoH1Pij8ySdcCVQIJ1LZaY2hw8LuWst+
HhnzEJjbHGuWUCU5j29nZ7Ue+nVLdZapP5LTiHKv53O5c0EgsdUeC//mOdkZoWRUk0sGsPSaAtw7
KEx67PizcumSxhlhQpYx4KRXJq8Ip5LSzOXszwWKFuHWnIlBwUh1HoefY/s4zBZphhMoDsoKN3if
09Ua4+8lrBL5Y3iKd4cGaKjWq1s3g8m+oj43rCcfknw/wPJn1Ko0b2kn+FuC/h4r1vD6ym4P3HNm
oKFUbLnzTczecfhmnLHMsJmyPCpYffr2yUSDxBCva1UWRDKEKW7qsdtAf3cXqJd/eKLyzq8bOYA6
cLgTDxoxEWu1/4BN2OOUkcW130tC27EPg+s7Vq4l3WsW735tiihWcoebeJMZBudBpDblJu05Yo6A
PqUG3jBc8SMfH+ktDctd7SqRSEd5Ro7QOsbNN2buPrckogUqZbbOOqs0gcah8Zx4RWt1GEwLtpmm
JNIigZSIEd9CyDX4bvqUb0rgdK1J0jMr+QXM7IHv96Qx44pcEiEs7a+sXViVnaQguBLDi+SVfM3a
ViN9Kxy7yfO91NmSVaL97DaMR2hn1j20E0/7Jptc0mD5TLxqskp9e6f+/SyX/TCuBQdua7+K7gQY
+zaPcYrJdkEeEQA2NcgZnVj6cegS029Mc1VtPzvaNRX1vO5tGzOKgP1ni+ZT1af0CAavdpC5YYDl
1BYZH75v0tHWcCR3jGKnOUvU37gqWYcSTq5GooYazKi7kYCKfxx1zAyYdcCyiI1vat3wflbvhAzW
FbFzLlHwSft6FXUPcAvtzl/GoZ9CcebsBHMYwRaA8lGu8dx3cNSkD+tjZSk5UdsFWsQZi+z9zpZO
ZPGaT4RISEB2whc9loYCJex0R5WQ1B+y56yGfFqGmpOV9V4i+C6V4I6KmeV/L+CttIXLgBAAsO3D
NZWYdc0jHuDAzZVky9G2iVVQ1ZYrAK2s0jR53SSOLaY7HMkIGk6aVTZKwE63CcorRiJCrvjYzuvF
JTZREhlVB2czwlrsRQLG+SbOvdiFKb03x8qp/ZNXvBZuCpaMcFBmvU8iWn9tVRbNjDQPEaTNwiJv
3Ukf/UojbIAsRe1lu9OBm2BeySCONS7uD8NTrTe6hKn4NEh/BKHj++S3DbWxY6HUHcOf9bRow4vp
0IykQEB5Ep2b0LAJkabssiUeNpo2UW+Y+tFVA+zVOLWt3TZBu9s5921ia/kBumXxCZZRnY/uJNs5
PvVM3lW2sOuFTQPiQx3gp3GuG4o0sNF/lU20chbJ7JKd/yekhuLTdVfths38NgpBw7r7WnDS7czG
Lc4uDNosQ8MZyJVCWPThhxc3/Bsm5cf4SkGCGVXqPzY9SMjDQEsD1lTo+UMBmbirL6xYHqIkGX8F
buWRD/iaayy2S5r7gYbQAcJ1zjrDGp/MwN3o+e+LneYaLgdpHVNTvbdfQwPgibIaLUfM9qs3vUK1
mz2sl/1TZHwsFYbI7/04yF795RUDN5mB1pgs6DqjrTv1PGxX9Mzs8SMGQDQz5ratnIJShhmGwqqj
+0j3ToMuD5kGO4tDA9v9EqnzLJsFs6JTYYA57hG+rHxPQ41jXf3EaC9jA3xWJYevWmzblD7RQ9/W
N4p7kMIdQQRPVe8uaJRm8n5+xs0aFysiqON3Vj/qd2Yticc58x0hk29WIUcK2FcLbiho8cdOA63H
o3EBgeg0Hk4LI8R6/rXjvZ3mWKiCuvxT4DlJ/A7xiilTskbkyTghK9BExxA7rtwr//oeMnYYUOVn
6uwEH/p3is/9vEQpUxtpSKH+CHS4RdpKq4x0DRBr4gupUJGsFzOYJtrQFIfYLOM55bH9AYMbymPP
PcYq4czdIrnf9EW5xRVnnkX7xdt5jtdkoe+j8/KlzU+QypaXY6tpDpJYwvMub6Aib3fZ9ejCr+yx
qU6VZRmIjernh2kORNn3I/q01esw2/9y5R1cOfD0JEsjhnDIaHWy9tKbV68cr07CG/ImTqqBP6D0
sgyUcoxXwzjgcBqgyDzxJjFvoehVi+hg+mDXZIeR7EZVxBaBbyoidgLGT27x1gVWIL3/FH+JPimo
c9NuCDNcmjaC2sLH1qsbR6nEGwhC1G6IiXdeO53m1LuL7IJSrvJkU3TcbsZb/HOHyq/wkCAXoqmc
VQWSSTmT1r2KvCdo1zJ+h8V4b2WVgeo1CgEd+lDzrhdJx57/VHxdlbwJpStMV7ZGLiSz6TiMXEnT
aw86Q8kRxMofvY3SIUZeBLEZBu1IKZ1QPGsUwKXKRBRc3K8t54hDzDUNortmx0lByw6QUqIZGF4d
cR2Ql6t5rrscX17Ho+dRyi3x5Ehj42lvUo+mJMK+IBwrNcA+wkagiqstOrzg0cLgx96HQUV25Hzt
4hfJYE/dQG7WLFtAIBrQjNK/B9MYFTIPgwQ6W6ZI6e1tqOzE4xvS9Vg/v3v0U8kbKTT0gxvLDLow
fY/1TqkdzkPXP9Xs63XO5v260Tkgfex37G1rdNGhoVV4hkl6dEwxg+UYk7KChiauuXKTuIV4B9Ad
2/bAPdJquQakLmiP1sc9HR9YpmKXQulNzBid0B5vzCQ3Hlrv4IXMd1dRiOX5Iluiou9fVY/trxoa
vRdBB0hQXcDyzQDkDk9fDx0vEMvPvi8McFHD6fGFYwEtYsdopgW7FQYDAGckTqfOkltFxHSktLX5
BHEpUtVDg/ubgW+ZIkvPcK9o78uFJ3QBvwEGqSJo31XZ/UcXBIxZho4+nwtzYaynEs3ngPQuyFUS
4J9kisFeReFEKprc7U7uRILqF8A+N2e09+CmQ05aQ87jYaMHsHae3fE99fsXdy7hDDIYspoZTPB+
KKTfzZ6Af0wgNfw6wEzjYTotkrHmvv/+bduFpm049mzX7lHzVBvVMpjuXNNJjoa+BFVfo+/zi0qQ
fcUoaHgktPc87RLawmJ5OPoWp6K3tXSw5I9RngemvcecWgvPI8lO3ZnR4sMabcysaS5Tss6RgHTx
5CTTY4WOtgh5hzeYCn7vlWn1ALnBbrpqNQhVbGqiZeLAq0P/5K16I4GhbRt5m1oS3M8araqkJMlP
YRx013TmdVHl5bv8aqJbXLHNdI/EB01EqV/SYWJKa/kl22rDj5IWozg4Tg+Kmr3DSWGzj5TFenDF
cLD1RA7R1mD/N5z2giuQ08ZxqUXAKsveK6dUMtIMeazd0Fyv389a5qxNqRqvycGNwSFDqKKrH/be
oqNEhZz/uULrpbGLMc2U0oGlZPcnw5GnXrDpfeQmL5mBvykUGEwx9YZDX1/WlXT/GPVBlc1LLLr8
tvxJazhb++pFFE3nUfO+UCKXgR8Rr/Rm4x51Xi+bCXB4TP1aqfGSURlobARLqIC/6OTRTCkqOpKD
UQrsMm0/xpZG8O8OBe76unKzsNNtKNhkgydKD6XD0DrPzLI5c3TFQkSIqyRilHKRtN0Bgdxy/1wg
qQtNlgMJSNl8vnYsbDIVHlTRlmo08+5CNDSWt8UgbyuAQixb0IwBWuHQNj4Ad9KtyJPDIAYzq3Hx
m2DhAtn4ZvtsvFqzWxx36AkBlz9mphGoCpeI6h1cAmRM644qMnQBE8GisaYxzDipD7WYt3+j/wSD
cw72XMEgJYToOqkGVXp2c1IvIK/Y2qXU08bbYDvW7xGFkalobgYC1htnB00pbx9LqDzjJM1B+ZNI
89IRQG41qdynyI1rXlZwPkoCLKiE624iInr2BMdwRUsL21Xpy/ohjLPpBYajP00LpdhYsyoD9mDo
8yLBM4mRFd34QWZo2kb4kJEQb67l93Hi+H5gr4WNkeAL8kQT1knqVP62ZhhzwoJmZH5W1IhikI5Z
US7hx9LsOTGnFuSKpzEu3Nz2FjoMbcH/SDe2tvNvQyHVhQjiGtWnNtZXVEfLqFTXOUUg399osu8A
gthsjey1RJsEiaEessxibXXKjkxLuW92mlR80trD+sL7LJoLswFIlY+ymiUhdsFYBD4Y6YMBl61w
PAPZu2xwX1Whor/1IcuVwu7JdvRz7Dfdex26YcJgUBxlVuDNWyn+KN5SLGASH6KXkwvlInGxfPpo
Grb0AFJlIwtisEpfGORd43ENE0yV7/wHuNi/4mU6jydDLqo5fBp4fFFcBQDQOnHwnVi7F5XHG06K
gNl4aLmBQtxp/0dHxhKPK0T5tD1d3dWZY/qTp4137gJa4+GgYgWf41Shav3fWP4chOtgVNXQdzc1
/O4vL4GVnHR8rTSHMpsn5eVrbeoJBRrBwaW4zEefuah32F70gzYzQBkr2+7ikuuO78hQiEqdIbfl
iEFtKSTVL/SftzECdpxqJl94Q+995jWhFKb6PjL0dbv5VJytAvHqWNfSdUkOi8uRByVZLhh52car
up9i6dB7xdhMRdsaWuPMg603S+eM0iW6LmESVA0uoJLObH7ALroR5P2Ltkad+lrQIgXUUNw2a7HA
bUgBvy1zDC0YkgzaP4+3UNwMKIZHoylGRElMl3aFLn4gXN3f1T/2dNmW3e8RcwOqaUbZpv1FTSTf
rSHiUVoEFHFCPJenS7I1WkM52i4iyDEiXSClqA0Yaq3MVehuBh2+kwt1bYaYpcjWi74/X+Zvz3jS
PQUEymLRcVIEhoCJ2j2AI3WMzbf4jaCjcM0+euZ1Pcmf017wDGCT/iV0DSIR3PftHMWX74I6VJM6
akKFZTx6y3xP6ccLjY9aJcWI4X6oXODIReyTBX0VVk98XwTbU4g+TPj4pWeo0hCQb0wUh6g/PQHj
f71VRmplCtXGX2IwKer3OshGDfuM6dIluKeHnujeauAMFJEKGCxLd/fszS6oIeD3RSuf7QbttHfQ
RkmZa2THno16QjgaqnWUxz3plANWtNJA4oNM5JSAzFXkL+NYBcUduYhX6CTntjf5lYKgBVzj1rm7
CgIGsuhS2VXHCRqPZKrQK5xGZRTRNU09hpPzzN+OupNxrLimqPEZUfdeioN5YrxdhcETYb+VYo/A
mYC0X8xcbyYmMe1BpNEEuC/G2tmt9MTwN8lirgNSb3v7bUWFUcPA/gdQ6zbS+Gp5qSp4WAaLUfuu
j9OE+gs2imvAyPdc6Psrh9P9New0G4nt4hvLhmBWPGiLUXQgBGJX23NGQAKUPxW/JcOFONtIrQ+f
XzyFE1G0+29kh3ijNiytVezEPuiKA4oYAWFt8HqHvX8BSHbPfR2r6Ih87AcSiWf6nlRBiEzhyqy1
FaxiOWGCx+6EZ/K/vzNIoEMaKOVnpjJLht0D/2EzkHKJ5EoE3kyVKoozr+SikKajY/TZOwbLxJOd
3C9uJLgkYP0+sJ3/3w9cyb5ezx6FB+nH7Gb+TY0AGNukzN0i2f3NEI+eaSJE/7Elg5rymKvP0zuJ
UEcYP0ZnB3n4URSNZV1P4IcGECKAVxwZm8rzfQDqXEmCigUd/Qj88MB06dlRlM5b/iX6NmmxsD4R
FoI+g08hpE9f3UoTzGMR7tN8sjN9fiN8dqOwMaQWpPIXO+MGrXnix497Jn4QQffLyYj/SjkddUWm
kEgJ+xS1rEGCZDhuNCQn7HM45RvhZPqzXI8ipVcw5vyyqyYLm65Tl1CmzZlsJHaXin0fiSKf5+nt
yIsVV+RGMmU7YdanaXdLoE5IolTXy7pAEez9/gGEhGtwNE0a93fjxp3ADYze/YiGtR0FMZl+e1LH
TClZRIG0UsObsj9luuNNSckz3fV9GCkyomPyemf1p+bkO+tnCi1b7xS+TRQYRGWc5ouOinpeFvna
czIpJV89dgB03gQIAcWwGxUyVkDMKTzwILknegne3gmP3SRRPQikcseKW1VrnksDrnXKVEMKfrs4
0N06t+ICeqzWiF5nynh7Fdnre2aglaa4gVoql5nSBnZi+4h8Z3diy3eHAR97ZeyvH5JlQZrAZnwY
ID55XdqEuBb0URQyPFbnMBau789x6RR7+k+IESDf8GFhTRXlep2UMgthnsCa5nHfD93rJp2KGvTM
v8awfD2yG+AZomiusuyR7uBz1dPyWwh7nTMi8WYTTfG0GegqS4RCJpoSq6nKatA5TSubPKHe3Np0
Rn4g1NLKLvlnHyKFJMiJg26C8Yfumo8ZR75VqhkuApcWKWlLY/b/6x4GiUnJdFd13YbOcc0n7fhW
IekskM/3yLteaOwFr73p9NW3Tqft2tfoz44rLePyuZu4zOY8wIUxgurQEvROiHlW+iysEmuyzcM4
RXc+fP6+uG0DB03os9onKFvYsa7DaHA2CEJ0sue7VUNqEtdIYnvhXi3uX/pH1uu4wUMLH192Xl55
R7kDRgwlW2ZjC0l5+NG6pQG0o878ADbYm7HH8A1gQLi6Dz5by5qu+ybnB8NTAJnX/n64OMbDlVbG
NKErwJLQW3oBjiFBgrnPKl7F2Dr28HllQrIDxir/5CQYGmobEnNF/0Y1HtJNrPRAFdugp0NENQ83
If9Kl75+r0yoQoHix9sGGXwfJqz6+nNFVWwS3TdiGRO5mzecMUOLeJ70GWdmjTPNBS25rB5W4++T
0Y0innKLUt36mdB3Cz3q/vYA/OhDkjoPmp9V1QSRSKtEntTL2fZxV1ZiHKAHJCb9KVfcF5lTiDTI
OjcPIHKE4HqSc/QLQ7giYZdbdM5sr8Ee84kCZFL4KrCbibnLjogBcTDLEJPS9+S8uzYYRC/BANvB
n1Df5qj4iOzXWUc7w2qPyloOXmJhuRXuPFYnhjBOGZX4mzut5xY/l/SHfX3rh+MajoKr1222iTwq
+b07GjXk7z/la/1HBO7ZTfvqiB8QxTBKUIvDEhIbkjgO+TXvtA+My1GeOT20jqL1fA8HSGm+fvCD
ihyDsicWGgN4MQE8QUQa3V+KnOgHhK0BEQSpYyYsU7LzT+X8lqWfrTO9yoSZ+22UAtUckrysqMHd
TC58H6+V/woWc7rhjQk2wiw2WTKdYmU8W3YeIz9XdXMN+3suM8U8UoDqIbjAxWCel0SZeTMVphI9
D+2feaemirAl1LvYGVC3j8SvTpSN8YZ5Hu9Z9HuOo7OypkJ2m3yAbgH/wep6MJ4qB5bF+LYmpOk3
IHfdEy6+Uz0O/OP7LwQfX1VjoPAsb6c56C+0O/Caqh4e/B/CK3X8BNVecNvoWfk91Mv87k2MnSYP
zRJXSGUKp0OOCDe8PjQAitKS80tRURpsN2DPVBz9wEUo487JL+Il6dmKsXvGOmfsPra2a/ubcC+t
NjDDhP0/sXv+SKo3l0Ge1voq3zCxpoqlRw9Hlt/WXFAgFBRxRMn/hq1ilm8ss+kMCaH7lMMtvqP4
pHhpS5YyWzUjhgM1SDdmMy3MLxsMuPyEufL9A7gyNTITvKU/rIZYkWIUyg3/cdsblrprghExN++B
tCU9MKc3AWn9jy2uIxQmNoBZsn1UH7UoziMwyDY/cRff/QDMpyimbj5MyVCKcftsOLgnpo1/z/2x
ykxcUWEoHPJVdZVt/LKBnoWje6cEu79LZaM4Eaidbfi5fHoM6l3ao1ZLVZeb6QuzRaAVYLfSrAt7
hLkTa7loElVJTs/sY/t6Fx8A/rJAgbjoUE1LpwHghEWhCUNg7pdiNCL/zngym7DOLAJlnqVyGVHW
tADDIazCt9cMOy0ZFKqzPsUOSnZjR0piTJdwSqZArbR9IltlHO68s14ANtVuJwFcrUdU9cN97ufl
HLwjMSrcEo8+LLil8mUOk48+WmpKM9p9TZFFjLD/pn7SzyVikgt7Nz8cu+C5KEnoN0QCUSA4so8v
HQQMf7Bxe+Dh06cBUK6eRwOxfECSHnbx8vSXtc4BaG3rdTb5ebmY3yZ4zpnuDj/QgOCV644t7JZ8
oZ1y4eCFx97wPouqDf3PLQZwCLPiAMmwBBzy5UQpV8NCfT23dQCZWjmPfeKkclR+tyn+YMMqzBOc
2bUDVgtqI+pdCUoIYXlEyC3A9OQGRTLXIK2Xh9lO8T0G3Hg3wajmZl7Owt5lI7Svb3T9QRmEcO8F
ohlNRJiNn7TwWuF64dVMPP4BxgNqXofOunKI870BKehHrrsSYvug/TryB6Z3jf7JF8nrB1ypY2iL
AXoWpz9N3jR5oGfBrFirvG7ABmq9/KxWmkJU1LYSM64xXt0C94FvqlkxBFYJmz5IW5/6xez1/PCB
dUbJHB/4gUlRq7WjJUUKS3dCeM6fUvl3lkAEVMG672oqkneaILHRcM7Vy6I3JofbuYqp8rU2N0w+
1uBif0L7vPku+n2FNa9XKsZ1LktyTbIiNlu35siO2etouafYouINFRo+Q60rjxsUowsA7PipY/fZ
o5Ap85HBjN5k3Srqyl+yFWy/Sikf1a1EOksT/ePHUkWPM9y9+1sdfBzo2EbjHvuMINnOB7HF6wra
bCi4f06p6FXNRuAXqKuP/FhK+DI/NyOw0L6CCrE1Sn0KXjZoZaJzxR3ckIAkDN5bfIit9ebqyAIC
NwYIBBA4XpAsNSaXr8669a+oqip1eHGLfxvDL10FWAUXV17Q0LdWLua+qtjHLdPPju2lrC9C2zID
cOeGnOxEH85F0GVwJGrhCAiHgd7RFaH9K2p70Q/k0CyTXXa3I/6quEdgUwCO5+9YcLhCZvyl2Cgs
vbCgu31X1ppuriSsvmx1HNuSLSn0tbfWMG0kGQKDyLzzY0VjUeFKeXew4u/M1mvj+hxXxfZtCbfc
PlQ1NxEdYL1CPuc2PZMrY300olG6Ho+Xal/wM9PVK2FdKlUTH/yAi1YPHSKBc4CPQpd9Aa8fgX1T
3QGKd8E16CXsEQaBJeBqWcO2DObUIShxzqlbasj1KDtXyPVpHh3lnUxh8afbZq1LwtjtJ+ukWaUI
NKU0dC8Chp6GAIMhhh/YMwksCxAevCayJ9M6byGazZsfPzbbHel+blqt3QHC4+uq936ssLvyO1vo
kXBbm4OMv5R1gMVUTpZmo/dcP1Hh4i7WYxFu89vvrDL2Mw7hM5fDf0My44hA0kjwlbTQRmfwzQKM
vYIxpml/eClk+NqSed9/7cqBu3nlWUZ1/i/nBcdEnoTqPM1MALuSjRGJkAzbD5VU+o7mzElbrRHQ
xNujRskfFxcFklwsxz+MG+LdOJqCr667lZQLmxTFLylvscgAIcK1EMb0TcFmexviD7bxhDFUpr9h
MPKOd5/nKtSyrGf7/XBkKre3lqkM6r46ogLm0a8NQ5YUirwvCuYcisImLaUN+x7fMu7AmR2NLHpm
pJJruCVZQJFEcPjG5Eb/Wrd/RVhknHKwF/uaaGhamgZ3PNDjL5ig2Pix1wYzCfMUL5YDq1o5wBBy
wgOsiUYW/ZbQlqvm+IFsUL+WhO1Z4dbhNfEoZ+YWsGmRxvv3exf3gRytcPCf38SjBIY1F+FpC77D
EhPTenvyc6GK5fFaMKjnznZW/L/i7cRxm9sD85Z5JwhT4O97dSEqMF2/kbSjTLJ2Qr0YS2DK376K
YAahXlKO+S8Z2eyTSNmbT9I9zH/ruikTDbZMSt1xCS3qBvGmpuCk5uilAirGBzYIn6lhdsPF0Pa9
dbEHl2+1bu5J8tfMGR/sLm+3KjwUSXyOR5WxzDzAaGF4wV3mWZmElfS7bwMjRD6UByfUTMrKT0Vw
aZQu3veqXFGMGbnGrdDExElZ6R64xBlCjLL60jv2djhxQP1sHN+JF/Yht8jPDvBt40cQaXdCCQ3d
FnqCy3BMJ2reRrxgok+girjGMzinmdViJ9bYKbvvhzAxP7KLF5UomMSs3t1oZIQiELLqdiag4I98
QFFqmL8ej8i6Scr/IUDaejW17aiIwG2vVuVBJRbKszgRmyP6ycn9tFsZwy9EJtOdShKderO+eA3F
CjDAvYrghvazl4pjmjAGXkf/xhU+7QfyOOkZEtlZhKLf92gVrM8MGb8/+rx/YZfdYDnZQdqVa4z3
ZZTp/qVTt8cSWlXgZqpkVUUN4kS4J9ng87u/wt0HtmyCrkc0sn9pom7eOklwnWCiSjq5iclp5915
KyF/kcafmHGuouZqMBot28FBDJnUUW/SluFk7SjYMh2lArmKCuAswlkbhUaYttZ6/CffkflMHdXV
uf+/bk491mVSfcgkMhabjjw3SlbULfbM3KVngxVeRHswSGriZlvUN6oFSMAei+Nm6CbPf77DV21L
a+Ud2BRdMcbBdkfk1ieazd7oA4cgm3ZNp1evpemMqkCFxoUqWop6pTUSa6T4utv+vILSLZmHI9iw
DHE/Z3QWR+KBn00aN5qihbsi6RLviSyc1a+65tFBTS5+c5f8aDdLr+O9EBOvQraAydZntVkiqQVK
b2GGxUruQ09wbzhP4AWeQKYietyTVThInDQ3kHRhsGjPFZXEQlfHQJ/9IKFySE+u59sLAAgUsAxA
bW/Hm5U4OntNautBL7YuyJLzKVl2ReAVr5oesCYyERgxMak/50kc9yQ9dW9BaGglttuFZC4Ce+nf
K2ToPZ3jxpSzlXVVmiJw+TnTphoml6VgqXSXA9Y3g5SVe+s5namipW/NSmkSFNKBFAsQlMbQIQkN
raup7O4L5yeAv3UcwwhteaiTKkHwFiSjtsUVlEocW9UVbw2MLT5AyredJqIMquQDP2Sm94l8WWBq
Nie+HReF+4LZXNljZIEFQgilzwwOhX0dY2gNX/58KnKx7pUOc0byS1H+hYdbnHF+EBxikObDVKrk
kAldIDD+enJz872fnLFf/3SKTa8O9JhlDSdq2arQgwzRMar9rKWwxf5DGQeUVKylypsAF8h3zP77
Dv8OP0sFUleGX7YIxxLTKo7aCzHwTUaPRRQtFqf5vh+b/GegosKHbZMSAdDKIaUKv46w++1fdod2
zBRGt1edQ0eFZilsLj3GHgRlu6c7M7k65rikwEFG1J14dHyldCpV4N3a51lBneLB50sxcIj9To1l
VDFG/jPC78S0J6FlV9ewaZ8XzNcLNmOrLDLCUP6j733uMEzpHYJqc9lZ/DyB65SEX4LdJkWskgFr
YzgJx1/6ULiBF6NFlQTDiFrZ7MKHNrjBW0KJbrUUZmE5Lr9TL4R3wO1CPcAmkJwz2v+UMRl18emH
L8UROO14oFSVuUkyUbnQe/bpj3kA2gpBqxPYp38BDrS90NNmfRZZ1YkuVAvhU/92llk7c2CHModr
3JNs9EumI+6w68Fx5ATTAwrMbSpw00tfjYdR/9ObqRiG19Y4ZIcnpE772czE2iiAmSglQn9ku/1z
xmmJmUNUlQPW6XfyaNSTytjgHKMQ29DOnrUFz2WrApXehVuigd5ZcldwhC38AtDsSpY+U58fghD9
l5eO0wvlPdd911//yir7nF6adXVXG853I7RiF7yTCKBeUzOJl+G66xo8izOuIS5kADOPqBKVxuPE
JdbFiTvoiwqZJfB6M04IwBVN5wmk2mtbZV6dJonwdhZnJJp3PWQlEDi7pYwpCpYrIII6e3NKW3wr
ReaPoMbDE1z9F0Rk3wyDXi6vdytK+gHqvam+nrrhU8xNDtHRQKDAxm61MHOXORCRDhfy8QgNgQwg
te4YdhPo0JCjv3Enu/zSNyzXRXzqmq6kkm1rTIg6SlqjW0+WBsP+aHfUMgif5puv4tinlFr3BFPq
y6Oaq16tqPxHGVfTnHrswZo0TbeuxHmDl9QSBencaD4FZurnPyQ8Hn1UJ2RXEUkYTRXUyUuuKOZa
KHrCAXxJ1GHqf0qRVnNTNdFN8ft4NjY+csGbRSA84vGR4PZuGDFgE8rgSefgks1XzEfvAurhbM1E
FIAOgD6xP6Jw5tvxpSMOwtAtwS7wJGHYY+6lIwjDMfk2RhTqksEM8gnn2qIu1+ywUYA98zQ7FRnS
BpevdiAV1HQOmhvfk+YElU/amiwc420jokT1LAbXGJPLrJcUGvZE5MThXVkNZfIsfAS08+NSWPMq
bgOn4fax8+AzJKjvjwdTVy6P6xOzukUpMpd7ZMGAVO83T4ETeGElk0yp6gH9N3XaD6M7wajinYDx
uduu5c3V0wDU94CVBwUOoAAMCR6W+2mlRx4ZlZB22TTywBUxS0/XSsuzOYs6fyrwAJGuOlvs0Ooa
a14IFQFXEGcZLtYt6ga6DMWlnMB5Ou0ZVvwMHrkQOm+ZZg+JUkThlJ/T+IpGlJ4A9AWCApCzh0J8
+cjKYNYtJr5wGc2/o49xrIVvTjXSKtFPxo6MAp96otGw0fOuzhjrYVfNFoGKL+aNcQd6hmUIFNAY
gWY6lBmWVw45iuAeKVOgHrZEblX10K7MfAJklIB9TR3S639G0vL8uAqmxwYgIjQZTCz+rIP2p3ZF
Z0bfxvFe9t2cpdHFMCDghTyovjMPoKSKhwTpTVfYuLfAXeI9q+7ivNVtpYF02dd/U3JWdsSUZlNY
HcgzdTdr/yPFDTYxDpafdAsEYm07TlbvZm18Y3lDNzVErWrwrA7/gJ9swhQl0Od/t0OeobmQ1djZ
fxzvTJMewKBosgTydihrYSjmhfCcWLUmCQCqfUd8j7WVTvMlAcYFvA41C4ASD7VhV7KNH4uW3K1/
drL3wEiod0N6YKK+dh0K5FNCIUorW9i9QhFIuB0P71Bb7hQZPlJiyYnvwhFmWriBjNGMnMLt+Xon
lI4RlT+ZRf4drbU2wKb4gGDJs0ekiocPk1igOcm4gm/Zo8YUOF0sLs3vYKl58K8R17MdX2/3YeIP
BCbUf8mcQGLklLskPhpSuWs242ztbeVHNKZHs+UAvHWNiib0Texs+f7oZGhLczJSuwRGPGVshKCo
lV1D/H5Afzpm653Hy19y1jQOttsTGqr88uLgMPx+xIUEHq/GjVSud0VoP2U6cUSj2/W0tzhMOVNP
e7S28yzOP1Pa0XYyiugPS+x8rfzA+uLSnTk//foUoAit/MTzlUDc25E7Lmls+6scydZWtWmZJxZz
nsOE1qNTLnRtpAzenNfNOuTRZI70oGrQ9D1b/5u3dwpvKjXuJK99Yd4gRnotvhSgEB/V2d0xlph2
W/Bq3jMa8aiV4yK66SP4T+XR1l26xOqUdnR80TfKdxt9V7xyV38IlhLrm+8lBgSb1wbDRre8WlCm
vmaXOGrDA8qrsFbmXlur8W5UCRtmt1atv5Famwmx7PhxQN4ub6ifJM38RLcjwTTW76BejFs3wJ6O
La6A59R6nJm63y3JAKDILh09mwdKkk7ofsoFJ5XWo4iUCvygD7zm0+JmKPqGdu+k/N+r2+tBSnl5
1Wq5UH/tGYXbWalqdnTA9KUOYi3Okk/r6tDWtzd60GnkiirMlz9WbPZg3FR9D3JRrFWtqt6B9XRQ
li0rikzGq3mBq7XaGqLKop2I8hz0pHWujoGmXtmAxUlCUVv4yMApzFoEKnyDt9eOJ18awWWYKOJy
TRotvH0jga0KkbsS5eKONQE1njBxvV3wrQZieAXMgDSDE6/49HteR/r3rbjgTBP2UKJGoa+WJQzx
2wkS62VpJjTpJ7+6PMrjwJEDWr1/crF6F4vCZT1pF2rCjiFhqfxDZwjzMuEQDth8JQM0YZg5RP3b
WrdocuqXu4xcxVb2xVeikhz9Aitor7EvQB4+vogk7X5MJ+/xnxUUtB9d2NFzbPC5hp29D4SPhu6k
gWmNSHJeerapxO+kvZjy5bqJDRL9Z1AdAOzvix5rNH5XbmhpzDnZvzW795cpczlj/mu/CidUs1zn
3CL95PtHiHvVKhFwrKEPaSDb8nmugG6AYKwnPzPX//F4ZhzEiL4tkaE2t1/Lm89RcDLs/51sXftH
BknBUEuj89P3pP000RcNs41i/zojbDRZiW3JS8psulrAXjGM1KiFo9ahzMH4WXDN7/xGuK4rh6rZ
beTqrlxRlOH+NWwBWFzvTgQfadaC1d+oxPOEHioZHeauMGTwpyEycLSqIZFySmDNayj50liVd1tU
DA+Y/k12fjo/GbHhWfcLspgbd1lZKR8Otx34i43/1kP/F57a877XLWx4ZJnnhxtCczXhW8Q6qkTU
/6vsFqK/jfKluzPE8pbzsezkTTvP/Iq3omiBcNc5tdk30NMYImjbU02Ld1FZ9peVEv3/6noDcn7E
62L6SEZvAkdfZIe3p5YIJtk2x8sVJoBwXyp6IN6odhdKNhUO77DPDcHy8Oyu9f8dCtOAryyastGE
Pyaq6S/nYb3psqUjlVtGv83ltQMma6+iYRDUAtlkBBPjwaqNU8eOXNyuFtlcL2lxA8u1m/Tsc06T
tkgL7QAuqV4DsskpcR1D8a1rzjTFQOuMP6bJ+yuTkTeG4HaC6yweb6fiV29OYGjQNuypaQVuQxWh
oHzCs4NzW9xEOSa24DcpAXgi4TfbkfdhF1/lL+Uh6XU+OLkVECtkdZmg8cM2wnwsNXnsUc+VAZq5
g4bTFlsE0MyAJcdfp9b5ESCswV9rrcl2Zzv4/gAESoxLLdOst+i3WMZbZ98scx6V3vu0bTYcIQvr
wcBl8CExGGbG2fypQRBr47ceQuElF2pqVKA25EI2zQRERGZrqgmO2hsshpSQFrt0M4vYTOn0opw+
EdF1q5CZjSWkLYQPAX2yeTajl3T3LTh1BBJypjmUv2puDUCRaaiAfUjihSq8ugAke1mUZ3248ZjS
KsvGU/x2GfwvPAl30TdmgsKOm95Vx/pGyg1+gkAUmZz4fY3a6A8ee1K8DTeurlKHLyHNHjnCp55u
s7uZoJJaVzqrd8g1CicK3SgxjFFgiBAS8jwXINOTh77dvSFswhHRvQlebFdkGEwEw/3f3Cnq8kqt
arCnoOdC9+ngRJkvWp3Z8/wwNY1NlAe0k71jiT0G685LOuxqBPeoovdInrMtOVnIe2jjs2dGqXDJ
m2rkqwzEOwPdEVMgSoAdyFoUm44f+xl6A9Qm7otPfFY/MZZ8aSin3qvGxU7RN7m/pWahOYhiGYN0
aaeBVtWTuXvKYnRC5Mdy2vRrKSxm+Y5x3xjiwYQl22I8rB353/Jh8Um3WcYBgrw0+20Avr96xkRW
NfA4zoeC6BzS82+9ZF/tdWcqh3aey8gDRISWgc2UPaiZIxLiW7zz1HJppSkn8vktDjJzhsDvKVCm
dd9pl9cDuhHyS29I1tmcge1PnoOQ4A60AtihfzlYA6OqnqXgeM9n3BwuIKyTfSgk3RzNM1yY4u6g
W0Fw2vep6dubyKdlKAbILypT7UMpnKXva0vf28qj+b4CMrJM04z+jFWfQEm4w19mZx+imU4SHsPR
1oB3Sqy7YEZEGx9hK3b3XLe9UHKvgmBW4hw2vEQYn8mBcqumWgQS/divzJ8ar284wRsMu0g+zGxH
nKZOob/aW86RVgz/+F66ptFdi7QYWXWKWCxVbW67BA+TELF6v2xia9sZWpBjjuiv9t10/UM7iOUS
SfG9Y2CtOZgPi+gfosGO3vcPiv4R3aMleoo0XCgxyVXuY5Jv8WStEsyCtDg++mBFjsf+ngr5LNKd
yclAy3ZuMDbNHKpEdOilzGB15qAe6gsRh9INod/+BmZvEg1oWly7PhOkluLhbnx84imDt9RoqFSc
iaW4S28wEDBEZ4/l+OmSG4aBUEFdwhDTZ4eY6cFpLx4eAZtS5tN2JkvA1sIwTw3N4FA0i9n1Oq/Z
kAt/qQZEFqjpguZ1oyaqHgTmxtUTPZCn2ylQaVtaXeWC7k/V6VSLA8PiHfZA8ZZRJcLioI3Inp7/
zqQU6pIIlGQ8HPOXLE5yfH2WR1Klc5I6E/e8G2IDdge6+N39n0ix/oAVBNp6kBD8w3LFDg0kwc/i
GBxrj3AlZpXotIjPoGi97lsptosgfl8ib7/bbkv7n/iVDuLhDi921fDkTn4ppVSprmhx6qiNRXzv
4XNHHMX+udwyloqWdHaY2/tz1hRQNfRI/II155Y6lpIMF2Z2JMk9pnFn4e8i+ghpvUyH6FrcREFh
frxgR9tzb9pAKJekV13cLLpPpEjgMLtUoKfa0YPNlET8JDuHXzeKxnQsgpvjQIV7g8Xx/xNs9i/A
rxB9FcFbHjW4BmOgImaNdbIZEzLEf3Cu26H530Ff3HzhI2ZIT7Wv2v59vCaCJJvXPovj32PPMLUR
c8q2CH+Wph0sZJ1neCZU4iJOnSAxs8yHcAqW8qPFLAw+CVl0E4XGKAVxUgldi8ZTDIHw8OxTv2r/
dC6EokoLei1v9KdSIPlQ/yQNT2pEWKAfeQZP9wI77EzvGjO4Nm6qINcqx883jGIMz9kTM8Vv4Fte
V5zxqH5+5mYvXsUEBfjNSiIq1Aw//O4EpJPyoZusho7vfIVVo8Huv8SJqdam0pfQPBkwHKcr+fop
NH4MURLamF2RTby+S5ABzhSbZuLUEUJT6jPLFBQbSX39Y6BzU7C1amWWWqe+cYvFdmcpGyk6ndcH
Nig+1wB2IIsAPW9/szD0oKAxs5sIvccL7ldMv+JOcrUX+/mCjqrg9oa728DTiUFkaItDyubL2NPf
MuLiimJo72eSnfCrM89As8wJ/qGTKonEG2UHFY/ufy3EWKcbo3WL7liK3fNvVkzYouz83CA+QQn/
iM3TnGROZnSpT0uiP5jlB1Oy+3UsZu3RaVXrebCxIGx5cLUWCIbXuaih4YcEE6NNVTEHBwbvp6CO
ltF8tnVGPHW2hmLMEsOHKB0Q76F/NmXYShHpgfWhFI8pUUsISih+t9wLO5Js1JQm8o7t2VLvWcMe
xQ0UOwtRFitltd7wWlALEVSlXq/DDDPgI44o4dG6yV/6W6tYpovwJ87BOpmFa6XjH80HwmzfB1h2
AC492PLKLue8NonPvJDaWBiFud65anPBjY7LjHZ16CKgk6oy78and7YbEnWoylhTDoYZDpkIMhhC
t2O13D5WJZT1tqyPSzhMYoropEcdA1bQk1PHPVLY25LYvLiLrdzbFdbOOF98p3Q1j5SlW99HdNlQ
snpRRobxAvMKuNxX5IdizWE1GMpR89V4ar3r4goYUKLT4NcaZgm5yQ8FoZKDo2SSuTIp+8ZlRLLo
9PaWbzu83gTMKvtBlNN+0Ipe4DgwkyL+vDGwKy/Yvc4r48jeK8N1bf0fg8gPolx8refwcq9BEwJK
iAsEQiREQRrb1m05eo9BtKyichOmFUmu3BsnK5MG0vjZDILZJMvox6HTkKc3FQH98fwDHnlZ9grC
kjmQK7CmBvUMnmtI2vZFBy5DW5adGkwfojLK0ZFD8/CzPaiShYPpd6lbq3p/XpTWKvYH9S0Ob6hK
0d1PcIpNXgp7DgU+pfIUL7v30LmLZ6XIWU0ahtCJNX4PuYalosFPxolUjYK91/aKodVyY9c8Ix5i
w1HZFnoHThX1ojprxpmHqZhfBFEh5kGicwfO7E0RcRafPEhSZ7VSP7edOHaBQRuGe6Y8HBbJdvr+
wm1JkH0FdEPTBYgwvb1MmFD9zV8mhMQSElL3SSCcvpQGWyuWnWsveddXE1dHpV6PsO5LD6UpExo0
q43IQnpDv6Ie7ImQHodkbaKLTwKgQPbqmWy/3XtdQ5f3Vw2hgIBT7roFPYJKIAD7UJOnx6XxvLXB
/R3tTHK+Ms13K99bPDhCEoVo/C4iRsYVUcgTs6qeYOY+fW2pFoTaRlkuxg08dcLmXAfXA1dTTVMn
1TpZcfj9/LMhdx1UnMBXJrVx9EpphSqUuLXCG71gJ81C2bc9bK1mWlS/4dPek6r54HzPvb/4PrBP
MwPUsGSMXU8yptpwmjafcxMPvJ4L7i3oKDWxeMNHHsLWmbdbNyBD0y3RWGzMZP+cdPHZhGlJYqnI
ozv6OVcFvcsEuUg0BtYALC1gUockQ+QdRlB6UvI3tt/mdbQIWeMvA1znELS11zw+y2eBR92RGTGX
Ipov2J/FV3dkWOv1hduhMXa5gFeo0ucKl2II9gYH1dZ/1FWByAkN20XtIYY0cAws3mT/U1pZ7Ojs
voPefr82KQ9LOWrkg28yyXAPZmOanfeFGfYJmWH5Z+gIDIh1SYFNi056e2aHITUZatmlx4kuzisB
xmOn9pCGHGYi57360XcngCxUoPGhfRchPF18KveJyKTKecs9OGsxJr1kXc+t6a9B3UOsnXpO7z/5
Au/CMSer1vjPuUqQcPbaCfeKP+dRPOpwH0P0uBlL6EyM16NKOBGVwkc4gq0ezj83oA1sFakGgIHa
3RfguRxrYBg6HmXXZ6HEu44GoFQtb7kJDbb/mLPq6E8U2aHcJBT2LG321pqoeSVUy/1f+/rE+6NX
4eI804yTYsXe6GlzYBQk0xMwNiQRhfU6idrLvFp5LtTrIKFQQDwjUxql+3QlktJQUwNqTTgUOmGq
1sJu8IPh/wZhI3IGNbjFANIq/6EzkPhcKsv1BERuN4ZuGaE5a4xFWz7U0VQ1RwF5DCT56nTtZQhr
YuKFaCj5DNrHgyY15FyTds8sZlPivT6M3sE8XfKSpv5eKBOyvJJLP/BK79WwpF/dHWYf2Q9NxPfp
bwGwYRlQOf7d7ImXoVWemdHGYsvsM3RyrluORD6OSUtM0CAMovmcwrOaFUUukxgVfXE9X1c2imPA
oRw0vr09SWJUi5x34WNhD8AnEjKrLaPDJKh/LYXoFzs9G3i83ecVlT9sYTqs+q84HBvyuupGaBTk
GUOVWSQ7hUx2aVDZxEKSqyUEZgd6/a25L7HqULAkb9Ufgjvc9OKBkRZjiM+OTvdhCTSPBV6X5pVo
DE4i5EvYbSPjY5OvLQNqUORf+L7qi2uGCTs7+IIY95o4OIFywb9zmMFjeJqiRXBIHK+3hUx8qt0Q
jdQvReE029vC+06mHEGA40RjLPm9FH4b4PusfOkSlpdTVnXu3DsFZ5+oYHybaJoELmorS/oxwjpK
M8dPZT394xvZe7/G4iMNYNiFZmFqgm1yaWY3pG3LT4bWFtTxgDGTXTAnXj1HJ1weZGMWurhpYnDc
kice6npiWF9728QrGiSsM/AIr8hIdNDTXlFlALSHMspYszKbZdNVoCjzQ+KqpLL8ZkqnuYuW4ysU
X7dQ3BB1Uunwh7TtqQurMEo39m8VgqbackEAqOm2RwaBfSib3uOLkBuw4UDoYNGiJyV1OWMkXkPe
2CfDQO81BSadJgNtCvGosNQrYGUrW7BGK4r4wT8O/wzhGaD+GCtWANhTJp5TZgqjB6XJ9+Fcz8Pf
Yt2qGwEuGzVk0Zv0X9vgsKMe3piP/nWefd7N53WQJmQrw6x6RqUqmfgOiUgnJSr857RlwW+rH2Mj
eh8unksmGgba0srJesZcYSq8r4tGulvpQhSAOje9G/MC5/UfjTogzRwQyzqe71BM2XHZ/XbmCheM
tHVzZo3Nt26zHMLhyTvYyNijdLAdg6KdWLttP7rPevsuSJHtKTiF1nQSX85f7r6yP4asgJECytBW
S3ZOTRtG/NaFIAeVbXDo9VGfBqH1c/FRpwiT9xY/3zCH+/i+vxGnPUeheEwscC6OqKTMUwFuENZa
qeZhPffZ7rWRH+Z3PDkFAFPEu4rdDGU1DFDNMCfTP2ZoAHeigovjbko6yGHju7alrIPGV1W/OE44
PRnER9i/lLI5cejZ9BKJe0UCgCUSw6/xewG4VP2AoYfUMPmgxWyY5VILpSVr+9HNDtgDxLY6/g24
hkl/PLu1xEqwXom6DGz7RZPVcUU78uT3iCFqKYRqLsLNUgqudwVkR3phmodXA+m0a5lpzRKP06Vd
P7W0FrOCm+MiRaJkk2ZrTcnKbCWhfgUMtJjm1q/ZjhfbHIr1J6pg5R1TiC51nXZfRjc+b3/5tiSa
IY2igpoZpCC2t2Fc53Dx0OJT/90o4a5l22ItHx7L9tbt5UBPG6WMmg5HXgY3KcfnR1sTBJ1c4DWm
dcOn6m3kQalcYrK7Sr2d/OLiL1T63YGjpqe5g6l2Qg5qsl8aVVYEh0boOTmeGVytD75iiVyYEVlW
Hyooin9vLBXO8UgrXplj1+t+HFikDZo+yRC04IVs99esfMmvz/7dU9ANQ8hdvvapkDZ5HKFNYmmf
8ss6b31IlAzTVYAOvgxkUf/0r4AGyt8FXxB7I67ZF3WulCWua1xY2ho5IX+eqwUTmWF05Pozd+o6
54IN5sImpOMQN9o1lMYq4w==
`pragma protect end_protected
