// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
A3RqwIwMWiPNGHVLLWNHhbls1nyu0fjgHSES8qYuqevPckXFMKZnFb5F30649KDHxFrVKUU+v1WK
ugkDzCUOzZYnge6YdEjiU+dhrJNj0FX6/EWLHWHMCS4Uj6mF5YjOZRfovphPRdmmDFQUak//HenL
ouIIkkEhGQQyKQPCRZbQcdURjtLYkf3qxVWGV6HV/KU1ZLy/ig06j8gYvYDFppfiEZ1VPGNaVk4m
3gp7XlUomhnW2MxSF2IDYeoNWvlwOaDaaKqXxMdROoJ2nQ4orjx+CsEmRyMNXlQX0aMj/JvvLhpA
tcxrIV9TGLngCOIP/oRhvbc0DGWIZCMo4dxm9Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
nBxGyTaz3gpTcgbHH/+VXmhpmvSl/BDOF2hZMP4X14AHiiCo0dc3yed+ERdsAkdtvWaZTqUx4x2X
C8oCKEyVOWUSk5Zp7E/zEjKDAaUt5RdLYGeCwayETxRk0EpWCpTCI/F488OX+kQHfsSAdAKEbWsF
2pOygvAyZC++qLU7UNjBpG/orpyVMY1UKDCf4fQ1En/ZZPgY+tqUMhyZtLhy/+uKr5Vm5u6AglMI
SMAkTkyV0bpREZB1PJqfhCuUmeUkFv/Crhyr28O/nEnXbD779onhInwCIn2tA4u8R0KWChmuwY4B
hPB9p3rM2enjHZ5mCdHPFL4QKSC1kNPWSISr76ngv52c6S5CITpWBLx1IHXrEgdW3JXThigN9sez
FaiUJvmH7VVJzViWRe505X1Nkr5PuPHRvnS8ers44DiML6TVcLIOz0phN7iCiVzqL9kQeJXe4ulT
qUZT8zDunTdkgupqZRGIw8lUcHa/OOgJZo45aURCH1i5G1C3iyzvzp4GU1AansX0UKfgqXHwOTQI
jsxMVTH1oMbhmUaDJhrh2zUVcbSmdxZ4wWrS/rwZ0EktkiSIVixiUnyrypfs3mqGUyEsFege1VgV
ZOg4ltVZpk3N2wECUs+W/9pnFCdhrhwRqA9fnXHoWegL9L41mTYhA0rayJvYNc+WitSgY3Zmpp/P
a1m7lITP7KupMvb7EctD8HOPCUiTAfPhfPJdlJFNhsuuwe4dHHcMtexYGAYblBN8lZHyOCOKjMOc
f09sKdvSCGttnoTNupJQnm5XGJjtHHjgKHn0et6l3/NlbAqnFUu2qmovuIhjgv3mb8QIzXHpcozY
d2hk5zJJwFXNR5Og7Fj7Y9mPjCEE22942F3x6y0dmLxiF1N8yXWxRkFS+K4X1elA+bl4hAfNWX70
66ewDFMOWFcxGaiyqgAYzn2C6ga7tFL7XIlPMOP1bP3DCqu0ejU/rvrfJJ2EVz564xnsWqQp1XTO
nqcs+v5Di45Kn9+JckIxEzbnaygQD4Oy20Mjh1qK30LSjVyyzGhcYdc5x6xoEFR3r7cn68PM/5Pq
CG6mcmYMqOBnB19ydIaswsyF1U7fgbogWYU5wSH42B27+F9/stXyfsX4YfCr0ePuZyyriC+5vQXl
nZhJVT7kVsb/LLro0iwOzbvOG2evZnATMvefV3EdCGr1CvLyppsumi5xPh54qvLCgMEPz+luomoV
LyIv6Cenddl65+UCWoU27Zr5fpaEA/I7SXg5t7f3gbHetywz4EYzE1W1bTdsXGyu0zG7PrKxxSCA
fyzMuyLM3UhG2wo9sqnPuh3Z9e77ujyNsyexAW2x4tkPRoxo6PAdb5p2MGGtrRGbNIemE7Bbcmr3
WYoVuvqpWQMsYpBYtU3TrcPLAX/atAf1Ov5UT+b4gM7dTNWWoTnhPY2QppmwAJuKogWPDJBKmfuR
7UasV65Kjy0xQSKY3izqs0FsXbAbcXwM/uSqkAa38M5Ndps5/3k+Y3S8pshGxmSZtIvq1xksc4Na
4+1w8HpvRnr9eAYI1uodATYc7p9Pg9fTIuFMvLs2OG4ctEHIb0AIakHApadJEB+9OaNlqgPuJkkj
AWZED1fEugFK1i8J/4LaLTPw3eLrdv8yP0H7e9TKuXg9hYtiCS8YmTjMgyUG41LgueSyhGJf/udx
FHPVoSHl5NRAbJNKP9pfzFdYK58GDWSTW6fq5JUXZMLrfChG9UbykMFCX61YIbrRrKBJfUHf+tHA
FhgcvuQdBwwDC6VAcFMyTGo3ET1B3K5PAALSQzNgzI87QGdcO5Rlzqitjb+WgcWNBFigMCSE68ev
t+fbZdZkJrFuQNS2cEJNt6XjIF+3hnFCJJxl971038cyuYXagD7DOK7Vgngt+qAC0ioIsKWjrDe0
zCh5MhiTkzmm/GHyP443l0hrmetQSsustTX+ywKNhZWVq1eTkD/3d+nX4OxbXJDthHZha78JLdUW
PEL9mgrIARCIkcyH6lKOruB4yy6fXLNnsszFwyCpzg9QsHFfseY9XZtzoNLVbT1g5u5JVkvihj1f
0+a3kZ1OGks19My6EJBl4Q782VfiogqIr3BKRHtU77BhPRbRmybd0qP/f3acZ2V4yxMcy7xyq0/6
2wXPEoq338X9G5avx+dcR9EniBSqGdSggOuyY5gT+85UMVRFBS3Tgn6UHNiIeShJVbqEsBaUcG10
GB04VXYRqJz+M3m6rRJt/0VWKorFOcWyhqsyXgjXT09eGNy7n8QcIMqP5+auJUVxjHj3qjzQieGY
NtND4JOOOOjdwpGkl9f8Vgiz9j/W05NEHjgaJ0cIVQE9+xU89NaqYSbvSJf5YTH2wqv79gL1Wd+n
DSxR3aQC2Oj5cBxMcKDFkzNn/EJLFSEOCTFEMQrgAJ9BwJARge7quoL2cYLjaNJJr+Tb7mYwO1dZ
Qw8M3CJTh1HZ93zodV1nORth4CWW4JBesOTkJW5LR7DsyiyJ4DKgJzs+r1kXxud4ZT7o+Ajo51wZ
trNVzVCEu5wZ3LW4U75Lbf2V3PJl/uwoYh8+j3GgGFpquqIqf8L254X//zdDoBle+olmGkM48YQj
aUgLWVmZKeAaU0Gk5cm8miAl+KMDWc0/IPTbyUBS6dC9oU1qSa40cWxPyTD4T7CBDO8dEcwtQ9iB
E5MAqTWA2oXhjzYU0z1QpP8eMaWRsjCbFYvxOCuC5revbGCHHXikpjINdOFbVccjUbG/tVThyieV
3QeosHwA/RonSfsVaEB9W2cvO/x0f7qsKKxTEHCImswuKapUPKUZzWxjzCyMfeDVrJgW1Rgo2q63
lGDEJnHBqrCwZTs0NMMXHMGfinRE37wEhTatPwLT82nKwwY9OjSXcfC4rWWVGuyiTT9Iq+yaqE6y
HTtsrKtS6bJommKf3oN/l8qOy2QnrBiWlUeV0Y91R9n2PD1L4tfWgYJPZVsugLSibHUigQfJqbGL
LWTVEmx3sV0m+qcmXxWvnID7LTmDiGJ+NHhA81e0UtTwerK4PJ8JMTqIAbnSkqRAa2kQDkEjgVGT
u+23R8BbIyklpyNGxfaftfnGAD8Cg0SRm425ttsHvEe7vUUKBwHsVSs4knYxYNuDQlh4E2eb52Z4
txlQIqiqRtFqL7rbCVTwiXZaX/eV2gBQMTAPgigYJBS1y0PxZBDXTMpb2vypU7fIe/d6jO8sBZiZ
s72fEXKiDQytOyFGW9jFWN3KGIWHTocZ3dNGJmr8eQhgXInREIDZFGYukcczSHmLA1J6bcweWOG3
u+hMSLZMaNsFTSd/CaVH+SxjwMNYaxf8MDB31KGKbOElCx5A8r1KTyqsgGREVM4g6ExPqf74ex5z
7DLu50aXt7Nho7vFUPJA9wI033ahoYjB8dXjKlps41nq7Vb0pSJo3cSPeCLWbbR+19NiaHyhipNH
nZgjyuMzHvwL71sxEMJqg5zcAsVHDKIJXCOW+Ya939rqf40BjXiDYXAhwsJMrfBEMeVMZz4jiAom
CkHPgeMuZNiu4N7rxlZ6RMfCbgRvdcLsQcOM6vfqPEsSTb63g6JL2rlpqtLjSVgo5VbIY10DPoY+
L6FYoJovo3Jdd7AXFNvTDjd0/4AGDwftPqcbuqHf5Tgpy0IjcUDmMUSOKB6hrFFeKH1CwcW+PsL+
fa2vltLk6TGEptQw9s81XN4jDsC7YG97bCbf+TB8l4DfPT3kIOeY1oqaUPBvwHxTHyR+doggJgog
L+Ymc07RJyaLVHdXsbqsILSnAPtZ0oqVS49PaSYqjPdVLSNoJJm3skUF53JnkkeUAe3O3uAMVxyh
JPMmzASZ6F7BL0FlBCJWKR21dz+AaOxbIZGKqZd5zHObx0vy1mBtR3V0rxlylds/sdAU1s+XDcxy
460xO0fQNOslj6G0lLLI5nHxtcU+t+j11PsvMkiJT7QbezTgszPouIGmJvoxD/yjIiFy68fTaScL
geQqCpZzNJBPYPU9PEXUi3R3WqkjNPopJgmOe/+PBijdaU6aYKIyqQ21zWVyhrcA1NsPVAON2D2T
fNyGKKLmksADg2fT4rYewgYeRNLYenYrrmg6pi9+7VN9WS0I2peKXwJ7Oy5QopZ1pC0Qs6DTtaPa
1RVd9nUAiftZR68NMG2hy3iKTs5rnBIe2nlzpJ5CkkuWVw3DYyqnH7TaBngJT0S9qTm6rqG7IRsl
LUtx/XAYhjf7Eqa/u92Lf6Rb5pT8tUaa+CM9caoOQbCYgKA9LGOq1oi0AI8vBrxx0csYEw7veQ6V
COvJxytA5cCqQy6MOrBduBTQCP4Y28l+jyC9rFARidgzqHpjCcdcmBUbwYsis2HIs+zsv+U3sUHD
Dsl6TG5KIY9PdfoER5UNHLG8PURJGWNbbSKj0c/Dhw7ZTNpcfchXlULHzZl6dhFheeCcJ+K/DxGe
OCYqu96wM5DD11/PO55tq7nlkAUdFoNk0UOCcqLwGldpAh1LwMKE/cmaCzFJLXKthbC3uLSaoK8i
OqKOyohnivgEB10DPhpH3DxWfkobpaOaUsffszl7k5uQ9nWH1dRmF2qveAxg/apULKs8KUYlYlo3
Ey0vZXapSgXmxIuPhKNky79Qjo6W5stcnzHApAiNxCxrpGqXgarH5hg74Z5CWwyVZyv0g2AmCZvR
polh5wz9FT/t/VR60E1qS3j63bETpvjngIVWK6MX0oLRjFVYZAbUFZd+0/SL+i8rE6h1Nc5rHijG
8X40xhGrkpVT7dBjpyWyn+CUkpgfssimesniDsCWyfzMSI/pebIipRn7GfqmuyGzKM9TCbKokWMl
K+BPW3Ox5X6kaFZHvC9JCe434VawC+KtvkkocvZqgm9ynMzQQJtHJd9b4zqDy6nbFqx4bKny7zHw
r8ocCCPbxM5L6iwptxnVDxlDrNiGIrRshvnkjqS0ORzP9Ns5k6PbDXXn/PFbVWyqs8/gcsE245pV
IY0ryG0siUlgbGFT+On9yixvP4W7flw9RojxUm+6PoPno2qSiwbRpXGL6iaJuOBYTOicfPbyw99v
E4nFAGOi/mI972E8q6uk/xnZUrYquibSD11+NpsRDOMoTN+E4HMLjn5HcZjKbpTK1EMBUpCPt8bT
bGsq107nI/JiYMVsU9Z51Ah5DoDT4a4LcvsijQ6i07hrrxhj4DM+KlRMJ3JvhaIfzrUgpj4n9ryE
B9iRhph6oc6fC/dzejIJ25kXiOjkiJgVyDHSz4peoQZoszepEPkw8n4iXZmErqdGqhinSxOfv9ZU
KNjHimo0ngVriMJhU6Vql0HnYi0CDvMLkXcKeXoGcMLvzFpChrZ3PewYZqSFOuwULupFuLD7C+MT
fE8vsaWGcUjHfINXG6BKrpIKvbtlLmzVMZW/BVJMFqRAHn68QVKynCE+INgXSzAWLZSWCuuEMptI
b0g04T0v1sfF4V4ySh8avR5+AHYFkY+Bm49QR9JbG17riqk8S1kMJjNJm7CLORorZCrWFWW5hIOx
qIwcBcvpoZZmrHY31LjQDnFSorTVU00n/uY9bdvp+NbR4gPKAh4OciLEPm7CZh0PvvvwJCvKUvtD
nW5iV6cSlsD7RTcPsRvW82xMf8C3ftDHMz4uQm6LKGmxQ5we8mCnP6gieqqHtaPhBOqH5ggWu+P0
R+60sewrmGsdZNltASHaV6EgM9t5TYb9qIDcihFivHf0uCfVzd9DxoIwal/d0Y9n4OEHgsOUEzyk
wIh1cmTkYuT+pREKQ2hyJ6woYPWnoRdi+N2o+7fQdzLO2xJQYcO3j5W5S/zo1Df9gOjiDsez0kHW
klnAbzkiuQFezUN9hUtnhFf2ksfs0v+ccLhHeKugw6+b1D81br85Fj+K2amANvutesx5HikLht8E
8P1z1h2bgPxrtO9a+vTk0ePMlCImjKhzOIWYhu3nMOq7XTAMNg7aBtJwHrw5ZGun10jaJC8SOgIT
6Cf8R1zlagV/ujZldpIT7kR1/Jk51sxbXGkbKen94Cmv95wVhXUdyAscL8wl2SQOCjIfJvhb/hc3
8nUWPAq2moI+h3p57JSWFFrKnPwaUImP46HTLaUc6QHr5U6ape3/Y36ZMB6zWcLTB9ccaH8gZRfj
IwDRQbAXwdMt6ZGpl+S5sMtXsEBQfHwAfRZvJ0GXmQoWV+9lBg9A3S9jsJl1uN6KL57QoAlxS3gH
n1yMVa4WgHRHqnoEdFa+V0ickPA5OWPpl1+WvRpsBVO1t32M3RAZ3K4hNhboHwzfDdm3OfeeXdxp
EfvIxivHOFtYqxXxaxO6w9yImORBLPcTDZVvagvJLpycB/ZdoxKgAkUHNto7OjQf8FeVDQxMuY8+
y3vnyhqThEtlc3Opj2Zax2bKvKz7k2kCgHTmQjbBN0q67xk7A3wr4V/XIYbsQRXmqoUzNb8H9odu
G693JeZEZ72vXu7VNsG0Bq/ZNC4COUTnUglk0Xmv6c4EtYSWDb8Hge8GErVKR8lDUo4sy4sSsJ7b
vrapRg2lacgIJV4Cv3AZVKWqMRVWLyJnDOXf4MGGOIQlKNU9hRAWDE9zutyOGtj1Wz4nLf4Y7JbX
PpOiFWgJyDCQSmXIkB0wH/2IDTDlAKmJfClOGH9iNZLhygOX3Di9mQVFvVzrErwNYB297MvmUk3X
d1p/p4ls0zqCTs4rSBx608SxJQikjxR9a5xSYMZRvS0ID4414cRfOllkikHnQYBfmWCiMYbSzy9K
t4qoRd5bkdQHe47A2ZNR/Uttkf9xBUYWS1U2m7iYFxNMHOifMu0F/FYFMXzZV6BaPVjbINB0aV86
UKw05A0mOWQ2Fo3Hh3Ci5XbJQXgMbfZK+SSVOX/lTIP5w3kQIo7gXf3X8uWVPtvR5af269NEG9hx
0D5Em43d+pw7jWWi+vaKrNIVvSMu66NXk7iovTGG8o3jToROZD6FV6yv+NOQD5RL0G5xJScGAjKd
Dh9h3+8XLFI/8s+V4/q7Cp/uhJGtXGbobrnGMjDtAsG7RSTnd6Gw3WLspa1hpZh3mYCuNV+5i6to
9JGSoOxl5ynwPk5YA9dhxqa2N3jbLLpagYe4Nh7srM8nZGOy2MShWpzsJJo2oLnJ/03BrQL9/hRN
lmP9o+WXa5ppHGHZj8S4yStivfSMRT1nvszErI8wPuwhQsFNngWXoCTHxXE+fC4ax/YmzzBoN7s1
etfoI2IRC/3GTfMkObetjAja4ASVM3tk7S28AC2fMFWkSknxG+F9aLL5fYRMFVRRlRom2BEJr/YU
5GX4VUj8kAWzIbxdoSKhfiEfI5xM63SaUzjoAas5x+MQM+ugCodmYJXtp0dXnkKhMP82xdDDAMZ2
Q0v7dt+s2Vsm4cGjA56vM+FTbrLxapellfCemRW3t8MTRowFOHXSzxbxaRmFOZzAWCisioOwNLoF
gQ0aHAftf6dEAv/Hi1RL6gYZKgeZ/vfc/WhGjXnF+RnuvDzcn8mhOwrQnIFDn79OcKQ99WHh8vQE
9nEQiUo2riPfW8S0o/aI+bkLo6XR4jIumhBjBS2sw5+vjAgl6QCG7JalUX4Vm0onTB99y1R+V2/b
07hqIq8FnmSjVWgII6lcvFX2OnEMO9FEUOfq9zbsAydFojxavNs7kQIXxzIrB9Fos6uzQ0f6MGbd
foDcUltdjVbPsPWV6UqPE2uEeaJHl7YZeuKmozgxXFBnLZWijs6F9IL3t/1Ieevh89j8xWk4gt2p
7JxuwvN64KxbD7BV/9Qcbj0CqOln6ERq8aqzzfNzG1EMJsyBE3sFPZEoqpjFuivdSTUQSsiV65bw
MD2+qx0Oc0O7TiFOjFczFsiZ8oHbQmLc2YuxZvNjnYPj3QRt4e1ShQK24SRWH+oaz/6iFEfFk7O7
3joWvj72mdL+yex/ugmjlVgNMORDTJaAU3HB7I1jShdCEOQiKNfegZ6gbnsHn3vIzcFT37Xr8oB2
X3oNJ7XvnRotEx1E9IN0E+w174idTujKJtfCU1L1/m9VtkVaxU8/5wj2pFvgHbIb7n/9Mr2LoqfF
zULManU8miXGErh4TxEv/FdmT52LcyjlANu8iKlmfhxC1EaXQ4pbiW5bhafeucwEOtoTtrrlDVfL
dswOu41Pmtg81OMH/b2xAtbXed71mPkgLx6hmqLP202OXjNLmvSMdeTtWvkvVYk/akprIlq6W12T
icoBMYZ4Q6663mxLAINDSkG8ZeT7woAuqZM130UqQm/GrTk/eDopRfvrdGtKbV+VSObyn2KtbE/F
KJaXQM823WDiK9tvang6GCcZgr7N40TPLIMEIdLUoib0tTpBT6cMWzAV6nlPIWMyXtWq3WjZsrcN
9IB6fPD+eNvktL8V5lx2424XNUNh2KRFwnAUY2aQKbiS9oRSXMTgtsJRHQCPXlMJA4GmHfJh0+ki
KEHzarMLTIthce4tfIY8uo88qEzQoLDFYxV0sNre1aq01Z34PhftSVixUpJ/4rdB8wmIu07zbKV4
6v8dA6aZ60NLf6n6tSlO3NZt8b2cnHWBMWJc+ADaEUK4ECWctH7iZnSe3AtiKXDSSdDYCPUQT8O0
4y0x/r4P4qxMcoa+/TGawuPTum88xrdrxR7cnY/dAh33ZVI+RsrpMeCEHkDT0tgW1D4OxBhCnykF
RG4hKQW8fsYg/T0uw6MlnTRG4xWhzYxq880kEhQzIVoEYDKySItSn+aMEr1kt4g29uwO4AIXlIn0
rYDyLASc/2zqB7ZFCcj9yAdvKlvAQgoyJ5csg8d8QaxEtoO3MJT17AnPl6Mj+VTZZJHkIoUVKkNT
OC95Xb/ecYj7UHs2q+EDQA89XR+q+kBcy8Llgn2wyCt28aKb9J+tEPE80X/9iOEuOgzfX4kRL9IQ
yJrd8kjHC7E8TQSkfps4DdD1wCDOeGfGM/UM+wkUJlBYiZ7mC8ER64cdzCgmF2FKFyjVYWzeJQq9
e541WPCHdjYI3dKwwcBfFnfq7IBd2U6U5E1cx26r3RO320e1TxXKTzonEWAhpE6vyG8t3fNs8O4o
iEWhTUKpAmGx4Sxo0Lc3qKm09VuckMrkD33r+BvZBK5EoTF3sJYhyQP7y3ECXvqgmP9pTf5gxePd
1lxbx/HwuaUcznfwVx3FLgrh6xkDd7h7TEc/kZ9S71IwBCV1AW5FnhMapCwmFxBp/UHxNb3cQuAi
J3QOEBMD1YYJyfphdJQfWGkNAoSrQIKkzAoilMdN/NTMZMsf78qFpIbtojpngZVEL837jvi2qz/o
VehAr6vcReoVTS18/Wjy51BNMGeWMoZKbH1dc8OmpUYa4XRXeWQ2bDvSOMNEF5hGFUZQ42LeiB1h
N0pERB/Fad4ZSDP5YqEfUTeOsE71YSKRIZijkaF0zNERwaN5FbDfsxCVvyl/s97JtlXAWSiTB1ue
kdWmoWC2hQS1rWyhDGpjXb15CDWAA0KiwhkVEWAH3VCDa6iGkLv9y9i0cFbniJ+QyocZaya7l2Bn
DkOIc2hhEN+d4rH83y4aonKjsTMQsU7j4X8heFb+CiKYY7fbrBSxF7UZKy5QR0UpHgYp9fYigshT
rpaJXsZFlpyqRa7l/GNwsgLazazUlwk+B2njwkw9Avc2z/PO4awJzUtnjkbaYfcJeWXrvkeyoI4D
jZD8T8Do1He3lxgO7DEvuswr/i3dH1O3kbWmUr2g0JBiRrDi0MWmhHz1C/ihzFdcdxvf2i6ziz7v
5/fRUeMCDTcQeRFhPJGa42mMjY7twOCFuwtOYZWEEESQ8zaebG02nj52LNUW0+L+tsmozmrzVKtw
Y5lTw68sBDRah71l3Jiy+CvE9UDPbug7EgyeFiJvvhiTiJSdeyvORH+3ciJuedLTvfkb5fyxnI7p
Mm0m6vJ0o6GV0g1JF3ouAITxAFr6ml9X2eJF7v7AYua59obih3x5OgFO5PD0SSgyppoSo8T6GmIc
Mbar2QQrFHmZL3OvfeoQEPq1sZmuQkNQX4+UiZv929Fzqfc6IoyIFjS4/p1wf3nVsPuVy0QWrKJd
pud4b9yestibn5OMo6WanXwZ0vS7AwkdITufq6KLLQRWwMbIbjISZWJkjV6SLA4ewu+s8/4cMpQx
wrypCnFwe2GouT9uGK5LWol6Zx1rYMlIPa6QVAe1GK6wdZyuXo/RrcH/q4Z5F2I6kpvIAfv9+M7y
UOtq7MCAIiudascU2DjK9KorwnJNVP7Epn6ZEhV8PNtWOqxS6BbSuC4b706eB49dK7JsxGWz8LTi
kznFpuiykh13TZsCClqNmj+xLBKQ29Gvq2VEEH1AP5XB2aRl5cSI3RcPqHr8tt/rtJs/q4Zd1dxW
EJ2ofRy9WXeLyEOAjrudA74PkJUjaM9Ivh41hMMpyj2GFYB03eIhegusD0/2SJuXwvlsjncqeeAu
6oZkrQ3cUSXgh8+wLfGMaE7/9KxdRWeDcSQoC3Aoqoch04Ytrqc3UGoYOdEe9InNgiNW0adXraaH
rePW26/B/FRpEqYD1IChqv/z24gbqktugkFwHRzMCL2jgqSbQQSczcgjti6c1jlJ19aGGQauny27
Ey94WQOf/R/siyLuFjGntXW/chjSBFDQVxm550Ab7yotsZTah+rt2Yi43Ts4WmFXBDZZjiHkjfRJ
1/e9jF/YQRbLc6RN+wRhkJgiCGJw3NWmvw3vYePDKB0bQd/NuGaXVeN+GJrzxkDeogeOSlNdFHiU
EP11V8gD0FVJTTJT7gaHCL49q1TrQGlDw6Pt4YjQF0pxToAnAkxBYDcLazHBgpg/HjUU8D7iUglp
Igx/fZGcREpksaEOUz3K81tVdoWcumTgw4mwdLHOjt4WEFXCdrCN19Gi1SYSFodFhyQCTzAsWMoU
maEQJqR3DG9xF0Tkd2kda+8iC7anx0fVbtUxofCMr1B0WKJzgGAhTA9S4fgtXMwYPLIjUtT/vWOP
nzMbHOKR1bUVr+ZKdZImHtgtD8SI7u25WyR4QaA5M3/JAJxQhpbM1Q/Wsi+wKYcrqxo5Ogmp5hgF
sPLzOgTs+MacbfD0i0d0ULh7e39QGL4uCZdw5DfMbZMWXac/ogFYHxl3qQ8tDvpM0G6JKRf6gpsx
QldTgGyZXE+l9287SFl8FXumdcL4Vy8QhEq8XH6MdnBuLsLZWDlVzfm39d94Yd1GVEeMaBPGDQDr
NkP/unR5dmmFbNKhnJh3vEN5QXRM5a+60MH41P0yB7gJEW6Jld4wvrqghOJYVL5tLGtjePuaLbyt
r9XWeMy2tqvJzQyRCxH+u09AZAvXI1BHoELdb8XGFXEAnyGxfTnj14FrW3fHvb5m/kueK2OaUnPZ
njzYrLqO+bzbg/53enuGLn/jnLuIRk0VXR0csw3hLCyMgT3XM//mOJ0r2U4MkWCvjCP9Cy5ySt7v
VS3BwgNmH+J8/H5pVrbA9ChtVObU6jYwPvy9qRyXVi7wc3deTYR7DCklFws0DJKrxmMhfIN0jAvh
4yQGLrBvXr/HEpmfQjweAam/KdmKMxWk1WHKMhvZcyOZEW917i3kM1lZ6whUkDjSNEoQuMPc+cUQ
mW9IuuPyeQbRY+r+F/HhVODGEfd9ceM90kcjPPg2JGW4k0XRWmrtx1L61mRL5okUEuoREdTGCzUh
LiXhcJAVjH6dvcz9Q3BSRziHef9vTTfCkFJZ36OZEZGaZWSuPlqQqzTiY2+p+cS0Zkksr+016svw
4ZK66uPSYUxKgoefF0ik+Mju+Yiw6h8SO7E5MtHw5rdPsVYW8AnswfRJGxciP11DlKhMViwKtV0T
1FHN77ry1ZihjkLP/YQ4HuPmjUijWj5vQn3dnIwFjLnbmETrX+wAXZsnkJiV91RdcnLgfERILAmx
QXU2heVesDYI6cnPwlV6yq5HzJ7QSGDFJeejywETm/80H5ZzrbzgnPhEZT4mibfJGV7gETDM4Rfw
VsSSAcU+x6TYeNWboCok6vt2L1Phk6gZGWwg3WdRvltQKhXX09fbWvTKtf8MgFzt+zMB6aNwKrY5
sNklvSnOn6XJBvaZNOOpERoXLwMtXkGVQ+aPQJgMk14SrAAGW9nhzSW1pyGIRW0zL4k+OzuLhk5L
l8hKqWZkBnLbsaofFOoTHSfnOAHauGogyuzKQyOjHl1fT02Q1uHFYd295QDDAG0IeZ1OxujoS48q
UnVxvyIYfQhxHBrcWwZgYdf0KI2zEgK2BkEt1agpbmnU/2aYtkzUb1WR1LPllUetk4sW6fBjwQuj
7aRV2hgIT1Xbz1wqUFRUXId1RAvvCsGpF0V1KGqdzfFlcVX+/JYq+p2VgQEHd/u7wLEwL5P8tGEC
fMkmF4cy6p/1ITKvjSDpI4xcUXoCeayCGsDGP5rUZlKv0xRqnBi6KuUZG5aE6RTcON+81irhO5UR
ABJDPpeVxBb+JfdWoGXneOpvP+8dpGtv1bIDNWbwoTIpTiEfQe774wLvhDoBLkHdweTVRgioP01y
AKnsXrrgnXnEEQ2TFqPOMfGv+ozdj0o5J2o+0nqa4zvorXed18lOsebme1xjCFgjHDzDanC/aoMV
ehTxszsyg5gqqmMpihN4qIkIDaU10nYXCD/girt4c///tUSNsPHpPbdDN0pxn24e7XbxDozHbGjh
A08gtnwchB0AH2wOVc6YeK7NKao6psC7FiH1hzjoQxDmdNiKtii5zOqOr8oKX3e0Wj7+j8MEtffK
Yg6pvlTorXN9qY7ED2o2W8t6l5xrbBOInfzBIW0AWBA5MR8v9i+qYZ5jP26ikMqph+byLnDJHVjg
kq1pZCr9HRE0rR3wHQB+ZKWOuXeDsqpBKzr7YisKL2xZ1DnTG0HitK2nv/TxmXfj1qsvKssWIy/9
sAsDE/cZb3jZdQlGGMApK1XyKv5M8X912vJ6S5+ZwW0+fxc0kRaUge6UhvbkvGu51/sCf8ZfF6Sb
ez5hFKB1VjA4Ya6Ek/PrA9BT+kGbudZMA9iukXmsVNf9TtFMZ/zSkLuFCI5rLh3bxM4SWRZaZz58
vWKGHdBEzsB5fMPhKGklFFIGzdcWDW4SgPLqg3fzwrsQQysJAjSibyfZM+TNecKgsRi4pHcFS2/i
rqIRVUH1pFAp33j38X3XwvZ4X3j+Tl2p0nFbY9f2DgJUwCbO11dJ3nPsDiXntCHl+qN8UPxvJ4So
0wYCoxlOIj7FicHb7AOEjsbuiRZe5Ss2rKN6seZPIsJn62cGC8L12G6VDdVqSDgH+8o2rGI/Mrar
oqXZNNVeSlwQE+UkYlUuVsbqezf5qKB7WnAG0LGxjiToeqHL37QOt//ZvXvpcZXAa4kEYWl8Fz19
KgmnDLxW0P6OiEf9VcZbFLbp9gRcwqrglKRDN80kdqW19brQm5Fyb16LyzkD1XrSpxjQKsjPP3n4
iJ7tji35xBjmDotbvVn+CL5+oDH7GVh+fktR+aM8oS2vvp2wSJ1BSS/XDDKTeBtpfYwz3vwIb01L
ZAFwdsqRX0mvX9hEkdlu1bGDsACIM3CIi2WaApSj1HLdlJtIIMmSeIw0ZhXUAVXTm/xiBQkA5Axl
I68Kuvad5/Ua7iDyEu+lEYTYlATAc3K1IGaeAKjZn+k7Ur88LoZo+MXKX2AejGWFb3d3RWrG+w2z
zHnEYxaWM5DtyFbOYWOoDXtw5XzMHnSOOdaSE+eeg1byTxb4xmAHiTh+Pi5XfQsz3Mxek8uMQ8JM
MycMIHRvR1pOCCA9Wz4HhLEeZIe2cjEnG/HhBBPSXBnMYfbgkybQ2jnM47rJrHfTTE3deBHzOAML
xvMJd9iTE7gRU80qokdNdmihfPas9vR7HkcQSVFBwJ9PTFndOQVcYxsA8TGHEvcB0pS1uPIwUXhS
MtCzWDfNCq0oLgU5IHxAths9W0GssgU/ffyGwXrLS9wszyoDMOKL1sPlKDxiNRDxHvgYJkRBLU7R
ATXAgnQrB6+LLgBxc/E5Sf+JMri5F94IXCP3jDW2DC+76XjNOjwTftkQPZ1+0AEoDNXnUvkdkstO
P4WMnTDS4SkkeEA4Gdlgq8H8t5iaprDyzEeN6ZH4XrTR+jmPPXzTKGJYnWbU7nUlFbb3WPMN/sME
cDYGUkKa39Mq6uSsgN4Sd4oxnhe2reeOPpmbc0V/G5QmRqhjoHUhvkhRMbRvLCDOz92KJiLnbgO9
wjWDtLgBuUZzABlo3quOVqXB+JpdoTj7lZzmp/xSxHUnBZ0zvZ3RcBODcMcLyWj2WA4WAmjEvHxo
cTUueSnHdfGDMgt6lFDepxJFHBngEo3n2pIfEmGOX/tIv6892/beE6e+rzAgfy/gSNVLFOZgWEHz
AXeCuPEDJzkSUmPH/1MWV/Qt+tS+tBTtO00o7mZWFTkF+zvgyd54i7IN5z+YWu4RNcOkq/t2rFfq
Vdz7jKg0f+ouci8HwTeV/u+HHhJhapgkLJmUuYBn91jKfk8AZSRXid3lFxHhVIe0Go553HzPJD0O
4lNT2eszQgHP6U7bJ1cfM8Ma0WDuAJTJ0H4iQVKuQZEDRLtHEToKScZxm2mZOzZ4gkD+N0mDPjGQ
Tw3PoqmnpaS6DaD+49QfAUmg+8oUIk6bFpiPu/gaGZEEHxGhuDMpfT3jPyZgrod3C+EP3thV1LIy
dfdWf7o9meER0ExYl8PCTF3QlCB+Ky592LjRks4TQN38iCALt9BDOGcK6w+t3GiJy5exDXbv5/fu
rMosDMP6/IYfIwD5Y/ipZEobjPW8T2y95N/1cqp0i8lH4jux6+eHWdCjSwzACwefx+zInbblrtRh
QAec9VwK17KUsos7tO8S0VCHl/c8GUHE4BtwZcLKVWat2jyQHDT+MNjpcXJcqGqT2OAE3MNtx250
VnAQQey006rcQOL3NLJx9LGmXk6//wkRzhR3cw7usXjwg8RsDNGGaU2aFMrUrC+imeBa+l9/EBq5
Q5We65Og725xmHl7r7fJTUvROTsOWoNkFoLxYOAtz2YUX28KxFV4cIkcb6gxfJRRu+OWQDNPSYuc
ZRuTYgiJfVJ7/DFE8cocVmnCp4IevQZhGwr7c3kESLBXdmZBaiqh6D9u9ZWMLo8HznkGk+VdN3HR
veDbKergJ5FUZF0+dLYc8qm63FbMMY1bE2Bd5fhuDj/UmVhU0VcmPJKupGM2Kb5qwD4aLnzdHE23
vFZhgUcF77MpuYtXmo4Ns/rOl2bIiEuCL1JTcavgWtQKySUFIeMNe8BMng9MpIxO1HotJewO1Gj9
uZMEiEaBgH98wdGck5zRmPanqhaUyMP1yBKL/13Ct0WmcgB9UhTnsWKb68AV6ENbikL35L+D+ve+
lHw+O41cJ+0PBp98KkOwtnGq+u8mci5PUj5CkXgBJER91HwzG6OrmNEoJlYa/VMwIMdqts5bDUpo
sovhPcbPFkhzwf5N2ywCs1IMAbiDDOeA38pTFplchBTMroeVsgEF9HAYglbrV81dL8OPLoAzwcju
1ZMPRlhRAPFUVoXrzO1zpg/5JbSjPnlqXfUMJqwPz9iVFrYNO/UwNunZAufBL3FLGQ+b/BsHTfSs
SK2lV8l+Mej7veaAYV5FAgSPGhv/Np+Fzlum8I4Ei+jyVKBU7mvuOplrk7KkVJtgA/aevfKqYidv
euzh5wUh0eTAWRYwutktkT2Cf27jf0zytS0GlgfZBnvcULsQJgoVcLfPjVssDNs5jXvRGAFe9IIQ
92tITbI41usLKMeLeV87I2ILb5rmd+9xqaCltoRvDYcia6XGtHZAgVKI2GFR0FfWJyDQYtsqJGNV
0qvDB1fBHHeXbyWJuq2RZ0Sf9erFEyiK3jgzrMHaEbzuD7aiPc9EuJBbqbCFo+2OyjayfwjTtkJZ
YJMA/vMzIi9ixG5wzysuN7F7bKcGFZBGNGbH7NKgZELZHUYZYRGGVUkdJJq33HuMwOXuNMivTJ8s
JKwByoumli7EDl/aOeWV4SoLVg44s4IDUEJVaCwiOezNbF7TCO0ch/VrWRVnmhG3aRjbD2T1C1K3
Jb5mA21wKd+rbRGbGrEdTIumomeRH077K6vetLnLbcHexxsqNLxKcUi81U7QAxWow9bX2wjx5LHu
a/n0QvRR2lfD9RAMNHgBE2PTGgkDD8VtXCS5U84Ys1rnG5q3L1rlbH7+DYFoLolmT+k944qumCa0
3eHPM9CZLRiw6U4H3Oudlo24YQNtiVa5qR4kUq1HlB06jD8Jqu9mHG0TSCbO7hLY9YNsgycbuR2r
KjsIfWK5W69vHWjQKTtZvX5tSFGkuW9Gctc+bu5RU71d78T285QVi/8a1KzC2OHC9cEETXFZouob
WfiqJh48I1v7uJzUexzyXn4DHZFI/IhYkA/PjxNvCwGd6YwbEJjgErEqTo4y+x0gJwD+7dNGVE34
2qwfw1Y2SB6N7CfzTFyKC4AwgrVHrM61TekbZbp9nP/YgKvNN6ZcRUXGVezRp705VjWYl/vzZ+aM
jCZqHISZ97tS0mF3RBMzn/AUKKIZO5eNUrETaIKNU3L9+7z9VklT84zdwYkA2ZhQGAh4YptwR670
nYvwRt+rHf8NhYSFdvTw4RciIhVeOUusOvCSXUaI9Ks6ujrJSxKTM1z72gHh5TZm3pBggaUUsV7d
XVY/SvUfr1OusLk4QmR9uhVFa+bFQvu47UwUoJSeDParZgNN64zD6sf5jsByNYdryJA02yC2qGqa
hE0KjQtPXQhtvKRbCUwhxG/mZgUotFL3yROtfiFnBEWnHW0vkpJ1sUBNNwwUCisCZfhLO1WaVEXP
ErAnAPEkfKmromkeRxE84gNo68mnfZaVgv9NneK1UPrv0m0m+QVBphdebSpOcfaMm1ajlBlJPxI+
F3F4melXI8ldhxOFSsoGwIwZ0/+ZwiiAH9F4HE07BtN7oQ3+1EFLwzjmSkyk6QoaArWDF3ER7BEI
EGNTnKHJt3Zg0UwGQwhxcjTlAXG7VnM01zof8keiYo5k84OeIXnPZPE5ZcrNtAaKYdBy+ayJVDl2
R6mMtDgW9c8Lq+thIPRB8QkCAXV9BPqEOWkQqyzLJNbppvB3tToZPlwD5hxgBREOxZkCaop6UGMn
x+7J6SSr6ClJhmV2rRQm0hwr7eTV26wpSWzj8Wyy47b1546qEZBJp9ANy21BxUZcKRuurZLf2WZ7
sC/6wFGl9bCLZGTVZJuR++7KCB+7tXlPEaRgZ/sWmC4bhMQPqzV/MVHbD/UZqV8xiYKH95PCixsN
ozf7y6WF1cvs0WVTdMDGISDsanvQZkn9SzE5RqFMZq/43Pi8ZYA1CAVoZzo8Ma/Jx4WgdZBPtpG4
kUWkTsxMNWIN4NTe0zxpS8X2PGW2LfqHIfRQnspbzJZW928ZzmWiooq9ioyjmNeDMElBXZWHW9xr
untBes3tnyw7c9X9zkHtPIMtPi7MBhJ1Oa7KcoUsPuMuThqsDicFizLrFJkomsCBQ/aQTMlYJ+IF
ThQyznq9O5Km+YjpVIvokkssBiu0UCamGQZXbxGZ6qlYCoITADk+eP4LU6htOEADHicGcbmEGzZV
LkiFUpY36uROHy39SaGvwiden/rS9MyiOMScwqeVzZf0xxnXObuQGSZP7Lzb6EuLPqFYIDX/y7RI
6WFz6eVx3GPPpIIdDOAN24NfLoXnyQRbzr3lgSbhByn+1vyoHiTs802bC7h1IL0BBiUprrsqJl4h
faYRMe7eQvFv35Vh7RM580saZPmUdGVd2nX3bu9FsizEplXE+FFRYcgJ0tDj28I5WXWRxFJgD6Co
6i+n5tFdWJj60W1fWJXIeDiM61sEZEVHEJRUJrFGRnP+XnbNG9I7VNLWOncueReYZuQPpThstuOt
e6GFHhACeE2V4jrGE4+Up//qFCx41K11uC09EmoEm7xlvd0VbhLELmq6/1PKyUzjg6xe4fcl83z9
+JwfglGUOyXAcga3KFcm6vr2bia+OP62ArImmMaPSiTN6ih70zvibaA6z0XgDGD+n3mBZ7W57irS
i7eVLPt0osCSukY/wjNDX7FkntzGvWvOiVOTgYFFGF5mtjyuAa3iDA29Qt1Xw9ByegcZNyTe8M5Z
p3uBlcn8ZM10va+mmfZDVuHMxXL8wf08hWg5tvbSK0NP6Hnh9flInKC8M3fTj8oG1oucb0cseKBY
+FGGOM6962BklnuMfQIB2EHABVy1vGRciAvrSGesJSXmNh674lsTYqRbkjZpYQxUOJ2xuw6Mdmzc
CzLEIVuShMBTPe+L8zKj3qBtf3D2R6WydlP0FFiUZUSmmCcGl3svVirEVpuwIPcSGNvhWkUGQ7sX
tDSC/iGwskOx3YDckQF6ow8+IDzqL9egW4OMGMOv0m5Kfvqb5NsZK9VU9rWdrmYH2mhEsyneXLyD
m+dN9l0ZZmciLLPXvX4U6OpAL2FYVHgo491GlB8O/mHMZIYBOKCeJB92MUzrGs5dOkIzRpITYaQZ
c1H/Q6DHCiAZdVX5w6Ig/RgW9utMA0a25r7OoieCB66xY78LzXvrDKq1YV3xf/0oLz+R5jBy4XkO
BaHRv4+rpahOTxXhrN7F5wy36SdSFH9wFhjBUiRrATLl6V695+X/CkQkJJ9EO5ozjBkbnUCEj+dC
FhkZLtGnSQNbe0nbqaa8nY3nG6YeR72qPNb1SMN0ietZgpAVRC7y1LmfvLgDxglSfPn2cDoFKrG0
6qSZN1fhZsh/vSH8h5mTRQ7/hqOSihDU9bMmxVprmnw04pViQ6W0XTKE/oMWZ8DotQYFblB5tqVS
PWHFWlqYJ4y4rddz5KLuYlKhbMHiWhsWGUWdjsIzVSNCm2e2twNSVQ4oKNwBfWcHm6fz27402RZW
aFNPrDQXA+m5a1Gf1IjcglTFtlHJFD//t/O9t94pnbDWlIuRFVFZTYbUeBhg82QQup5HC4awzTwA
MzY7ubvBnE7BJmwpKFw6isuH5IN595lYyvb/JbnrHyfgqbbZ/D0U8nW7djljXVwyBiR/5cMnG9Gz
7KPJ8TFfbfITo3ufPkOdP1aVHhbUljPVAJa8HAurG1fqCSCpsVOgx+dIOe5dTEZKyT0A4VYiLvOT
EfL1LvRtV6QrXKHdjBtvF7+ky0g3nbaG8UPPn7IfHNtqVMl7/8cLz+/FXsuy7LBzZ+4Sk2eftSwB
3qoiH2DGh35hS8hKby5cgHqJF7QB4rsRRRxlMxrERzDBWIn9sNPWm1AqjuXV5aBTfDmUjTS/U/UJ
E1Y9e8q4JCjVlHQbCbHOxZCWPUBD58KDZINgLYspF0Eg7tq+2d3/h7gerSNwLv8Vbri4T0GaF6LK
pzdV4znSWs72j1nDQgZq9XeGI6I/5xB6ZxVfVdObqnJUOAOq2VbjMlbbfZI1fmNL/atU6Zzu9uyH
7KvXd+J6a6WgQL7JPr55kyewTpTtcheBQo1cAOEkpT6PGrUXHVfBeI+rL/XtAwOHD3GichlkcUG2
1gAzbVQwb8D6razoxcbWrJpl02uSURNBIsPXFAP6fvYOgqepNqXTc4+s9oNqmSRgNej8X1a4VN/f
Jn9SDCH7uL+wi2CjfkRsOh/jFqK1zeux24VoWgqW3vRyZUlgjhYOEEvnl4fTC0EpzuOwQ+2V3PBn
2Dza2PK39nHjAr7Mg5hQzzK4JiNKAbMPzvQgKLJnqGehkx4WScWKgKPZsXvo95m8tb8lK4hpvzLU
nrAQ/h9bU/0SBYjWzatl1gsJQcScaPjFtpiVtX4u4hn/WRV3KSjbqyOLvShgd10QokN6zBLWzJGv
TAW0TD5fGxATFuv9+TJGVniBDH9d6zfJOpDYCz1t5ORNIzy5CK1P0PXaguP/DpzsINA0Ev75PFDc
mFvuNEu4KDsNRFvbHBmDzscjFyETf4KQ1Q74wvHcYck3zEGiFk/2juLX01fYA3dPDhsNIguisy8v
N+fxf92pbsP1mANfJcVDQRBWPxb3jZYkn3uNFwioTzCESoeodMFy1Des8jOE7gK3JCd0HAQz6X9I
hhWwgjX7Kb0e604ntJn9UyDlyIYwOcPuOiy28ygOlg5lSxlnRxIXGIR7fLnZxzOGGQvApvArN6ku
rdkX7Uq3cbVnTvkwLCGSo8SyyTK2jc7Gniip1lJFL2zB3WbXKOTZybxGlIz/MWFIIcVwsDZVJ2dm
yHh/J9Hn+DqmcdVj+XmLNZzJh+liGw2r6RWHJlgBqOEoJGe/DW2FMhsAUNWdZz+eTABJbVbStS/8
xSufpI7QqdyAH/vvYeNac1f1AQvqK9zs8TFCK4afik4DZM+f9fW6i9dQW2siD+4Ja/r8Gs0Vv+1B
3l1u3EhZ4/u07UypklbHqDbmEJTf9fT/VeXdfq7+AeN7KyWA85p7z/ovFMZwjl9uZ+o4TDLOHYzk
LjKwiyw1At57ST79Mx79ihbDTx5bC3bqxJKQSrei/Irm8Bdt3zP247934x0J++p1Bng1VfQJTgIU
A/Isx8goQNmMNmJ4nwdZFFkUknLo32cDkaINMQBiWQ9/WscMwkWgQVeycaECx3NDwZU3gza5Pq+8
rio4BSloKesbR2Y2oQkRVyn/iHjCOUhYZ5FjXhzCssohcesv9VpC2x0fBds5tOEcxkCtbwGyGyLd
DFSFl3lYIcgR4t6hJzJCO9g6Mu0XVjOhGD3Pl2uG2yF/ZCz1YJrnikBRiCwF0CiDgD6mXaTN+J2U
ShzrITF9j9U57TTHlfAfvTThsGkP5GUCGKirEj/wowheXgYJOfjACKcbc4Ss7aSrWaIR+agSo5xm
B4ERyja1650JMtfyr0KKRqxCQF/JSdTGeo6rHHl5Jk4bKLc7Twu3aztFyqQXXGvBgvTsqpNzREmR
s9GUiJ6VWlu9l3vfExIA074PK7uw+j2Y0ng+HRjO9ywgFHI+CiAKspAbT9/2BhZPjlC7Map171hg
8cQ14l8Fh4VWgm5Rje+QrQ1OXZlANBmuVNUOVA13h5jGeVu2/L4ACPDkuG52/Ivp2shqxRHkC01V
06OlBhM/MU0ClQbOs5F1ES3f850EYXkU8TIm44W6Th1zj2fWkNn787nc39TlKDkW71wqbwmRm/jC
DN+Pc+8Nku5Rhs72ufMpaYEI0rfN3dG5yv9n7fLYahxpuU10EcXzPLv1IyVD34B63JQJ7QLL7+OS
Q4f7mAcAbpXiJvUUMPD65idUMbuLaVjrwhG95qRIq82Hl/AAFiFUYc/LT+3TDBJWAiIbgtndLWCx
TiPhhyu1UycR2bDzGK/h6KGrRFBxHpRlGY9e7r80LPH3nfpdwgcyZejTjP7xk8gp8hMeResjz4jc
dAOSeoVVLusxLJokoz4nBvx8amNxdwPAhjW3F8I/UTlP90aGTUcbYum4OjFYN5omZQIhOw7xKUDj
5oXuQn+BUZApII31wNo9TWnu6pJ710V0uZym7vRXrObZD5CTXgoDZoSbk12ZlnX+K732oXSYgNuQ
M/qc0/TIZFUUyBoeXYeXQZ7ZKloyt7U/g4mZo+YmykWaUVAgxEd6DoY912cgd3LVO0q7iYp8Ih1i
BWd3bEsY7JveTpIUi8zqXCe0nWgqw/czGQKBjmq93usO+ARhJNriUkgJ9AhMy6Ut4hyPAgW7UF6H
kA1YSqThUIGHFVtdznKwyQZQEchEFSQOHXDWo2l/yeAD4ObH40B3ltLTNn2kkDbpqywLMSGA2JRM
k1KWw5tfoBwXVr9xgPdYDMZX/9QVG+iL215iJbGXYqzDrFK/EiJsKHxMDCGJJWRUsHh2i6Rb1yrb
GEwO8P1t8iMy3fgBBeeOhC6nF4qZ0LwHmuHgSyBWp0zocTGRzQElVxwTG9fd1rrlTNIXLhkzW0Z9
24DWqpL5QI++wzKK+Gg5635PWeJRkuLOtKzFLfFTfSZ3sQtkU/H7WFuHTqT0N+xZGhrBsX3F+aXo
eW7GrExMciFwjakmtxStdSX65yy+ihCCGos5+Z1x4azrweE9Lrjbmeytxa0EgkYc/I3Eibj/10dJ
I9kOxvqpYA5JdZc2i9EzJFk7aN1KiIM7cw6TD48WD0ZMpSmSWLpAUtxT6LjiBqMol5I9PqCuifz3
0rdY1MZ2gt9mmRz3w+741EakqOnHRAR9/5k14r9annzDoxnG9jZLydOk11RA2uasVhD4G0muk0hr
OXFmrrqh1bhXGeBu6ye+CH97qdUpZNTYh54vrSKp0Vvfn5hbBO/2inkjWmPhyaQKpInM9pP27tqF
SyfHRPXZt0hx2ZEkJXrlzS0GWnLoCqOQVq1gri9O99Le2TrYbLKp3/AWccbuI4LmyI521onv0Dbc
Cp3qwRVxA6PSTudVhN3eZjm2cZ79PZimptDmm6TQGKakEqw3IaJMTo5KwwaE7VUBrBJEE6hKUnmA
jn6ZWYZ7lkuhbyGn8Oesjn/H+JeRpGki8pVko02vvHttPap9dWKEk7jlNkrdIUOZVyv+m+vi3txX
a8iys4+8qWoSz4+ophSWKbWFg/pdRuWaCfz/k1msat3ZliYGeQEXdVUhM33SJ2FXd8PWEFztu3GY
ItfdtCgNZfDu1AmGIxJEVltkiJRiZLXsf04twAw9Yz7IzaisLP9I42mHghoJpFW+GQpZHfzSGKtT
dRF42zzFF+jhgD+6GEIplDMSYA2aMjlTLN8bSAiDxAVZrzRPuV2zxOAzGx8pWId+yDZzlob97vjy
Twki4uEBc1y/J7/mDsm2NwyRHicUtGJg3tu6APAi70E8g4gwGUUxTAabX7yZudaNZo8wfsz7sCz5
EVHE09aadmq8MnMfQCqsKnd8gx21f10X115VTeD4ERO3ddLK/Ecx5kM546HhphdORxtN1uL+Mnv7
1/HEQWZTw6jGQS+jEjtxdoZZcGyz1JDKY8xyWBPSjPv/CmRrOrEVWsYT8nmc5baXvbLPFk9T3eq+
4a4ojKmuKzcGEXmlXDwXTOnd88Y76XBxE6K8B6D49wy4s6t04jLHYZwdT8pfboDKXmTV1P5wiZNo
PwL1BuUjXs5IXVtO8T8J4ymqRXDU01Ykxl79sPpBbZD3Vb8kzUowdV7WbgsNcWT0tuLQqPrOXMDw
cr2hgyMfUoznmYuNIiy028wCJRcmD5tMjrS+9q7Git6WSyqvj4beKGFr/4pefZRMo/4F4j2Xh+hU
4mSVPh0x3TvwRZgTUxOqQlZQ41K+qSmP1C/p4X6JTkg80JP+b31QOxD2O+gL2z23hP+1AS5KFxY7
c6NDvYohMaLPsAKfp2P5gBhYIqMWUgE+MNPPDiv5iL+Md0ARp0zr8mG+FLtjKykNoVAY48IpxXGe
V1KRKSj28CxhzJk6w4BWI92s8PAwl4KLvSsU5K2gT8iW/VNuA3+A6YFRpkMv4fs6
`pragma protect end_protected
