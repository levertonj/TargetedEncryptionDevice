// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1.1
// ALTERA_TIMESTAMP:Tue Jan 20 08:33:55 PST 2015
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lds9tbIE+gm3bf0Ww0GYdGc52cQVmls+hlI8ZMZre2aNTYGuvHftiIWTX8RP1j8X
f/ajPvpE2MEdTLN04bLcUVz5misNDQ5r1EWlJ9/HhKcsfNdirC+vkM9QlSQ2Foji
BzKOPJR7oenrVUPKUrd7THM53+PU/BW/o5r6KM/TVvM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17584)
6cCqlJ21YqP6mgVqLe16uqz1blmXJzpCdRl4Fq4T5pdZUEEAkSx49KEav/C+cPsj
EQ2N5hiyHGPME/th5oprOOCgwTuDG+PJY7qTF4joxEGL+uHfW43txloJWB3sCDhe
CwptrcMNSUEpRnzGEVRHMSzmVlSu8dZGhDRKpA8YWAGKiuhA2KKRj57dIbuT3+kd
rpPny3zG/Kk8/YA2jf09ddRw6pN+vAfYo3qWC/oNK7qqvz/nEqwcvK3Heari5X92
2Jne6GY5ed7nKOkmS2A2FvOZkTpkoayw7c1EJSX23HtpnS79S5RekNpdpKjsRL3u
oTz00JikV3oAnihJEshNTRgl0Vx1Y658YRsEiF8FCSOFLmDaMhgRP9fpbKv++Csx
5MpqA8j2Pz/+NDif4zygbhG5IzelNMR69ZPibb1I5Scdkwnz3T0+F97ah5p00CL8
9S/+DQe7RURLKZyWJhtvjp7IfcNF+QiPBif6p2pHrchdwzLwrHoJDOLN1Bsq0Pb0
9PLOnfl/WNdtLgxe6XIGrXo7vjImw99LKrCCJLGD7D5pAcPxIPd4EX3/ogouSKFo
X7ZuxzPaUzlCiNUVwVxEnBlFCDj9rfA8CyqJ+boVN1gxB3o7ao2MTeXGAqjSbkNZ
n4mHNuDCTc8B9pbHFosI/veItF5nuM42rO84MxM4C463mzfQS0m1mkDz0mRojS4L
VVIJJIPe22Ikvn2KofvkgOYW6SYjbrxFYk6kUlWdW1tD9e8EPZ0Pxr1Qe/6RlPjv
SOpkMKxQeDFIxzxbK/bvLQczoFoFDXWzLZnEvPehLgMS8mInd6OE8WQmchqdQMPy
X8xC1v081YOun2AwpU8uILn5mJlFnSyRceGwiWjgyoG2kpAx8jXCPacblNpx+BAH
fYI+JewqJgSPcvejZoBFnH6IVHlbIPJO68lFfw20FCOrbutZm7UPo1/3f8Oz4fXx
PgCtZaCVidtJFOr6RMr1jkkWNluy0THVdNAjlmoQ8oaNF/usF3C/ZlHpH/WG7auI
l3wvuZ79Palm/Wi/bmtIdDYBtJY4WPOtsl2zHZgR57hIPpl6MZCTGtqUrA+2G2pK
ULmyhR1w0FCI7HpejyTFacA0M/6gQ7Qsjc9Buw+J4bvCe41JDK3eo107sZPhF80Y
U8MXmQAN5FMm5OZtuCLmhwZ18nR1A9uDgGnbeI7ApqmErj1IgwsNlm2/QI9uf6hS
KoS9GJsqUqfmmoF2rftYmeWNXnP2PL+iZ/mBoT1EYWZJqsfsYZAL7191KJuBkeh/
w/UczxFBP6UsfRbCeewfXblJ0lEPSg7paAKakqVaqsFvrXdlJMY/XdJ78sbBs3b2
50CAQ7dUwsqau0C+IUCn9jpsN3SyL6hKIbNbZiIgxjgeLrI/dfT0/MtNH1GhVueR
11W06nfH8hSQMoNcUKHke6gyinkhLm7CtjFQvicEOEfuzRO7KtElwg6pQ5wpQlXm
J/9o/lTAlJS7e1q2tORy6PjP5NdhIQA3lkozXHLbj7BTon93sHxfaqJ9hAjoD5XD
zRMvLwCv70hksAsDOEnKVr05CSGnP7nyQDkIubry7jP78X+LXwgT3N1j7PPhbq/w
MNt8f87s6whX9KFNozji0dTLmXpx2aPejxe0iYFJkj9Cl7w1qLMo8ICifhvMJmH+
1yzGWsp1lNciIRJN2noTg0oiaieNBZzwjyudAeTEEEA6/SBasKo4x1/HZn6WTqDP
X3CVWWxLlF6Vn3XCYrYvO0k5d9UrDUFxy6sRX4q3BlYGU3TgtmNoxGx8W537P81B
bJpan1Q7hT365UWrJSEWqFJs0tP8G88JaM1zjSfdnwVWc1TLoqSa5JWsICWeapHr
RvheNxB8RnGaybAl3hk6qvm8TYu2qTF5ghacz3ERgmTAKnwMkuGQIEeuDnkY5EID
9m68qypsuhUAYSjltjdin4Ig8lQHZqYvLYh5C2rytziJCU5KjxJ1o7MS2Hir7UkD
x2OdPeUXEX91A/mePhFWzXYM5cMr3uNLBLCdElFRByCa5hVT64wip1GKP/4QEXq7
uS7YgHtqx6KXnEEjiq+ti5/nxvDrZ3aPmtAyA2NDF8Txw0X+oO2IpcysXDmQ55BU
3HNnVyC//gSTENZshLJDA6ZxtYeVg4GxtwAIQwJltFN86DqRIuCmY22cSsP7ySlb
aSJ+3EarzGJx+g1clWg13Em4P3/YoGJtGDbKiASehEcYAmRhXY3aNUJ7lShCSQsg
66q06Xu6dwO+uIzPZ1M84laME0jxsrQtreh6TzRTV2EqytQH4kEgboPN8K7nUzbt
UU7P+SkQAN77nojhXioNkehRUUsPoFwcAzUM1Gf08PUF9iNSjbIkhXvdgpMAxYaq
92yuYKRv6n5OgzdGiwVXATRaJoHtmQDU3AUNw9IS/IWR9Eea0dgEECTyN/uppKHt
xebUIGHdzgfcnGGK5aD9m/6m54NjnLp4PW7m+UffsGz5AVTd41RwoDTK7/jCsKZP
0PdJKhJ0bwCWyGpABUAUJyNQcAOHhM2zxppsgBb32LgfBFFRuT3bPgAhviO839/p
TcIB83IT+X5bl4Fr/QtIt0Vvckqrv0rLux42uXRFyaHqxZlhUqSV1YU4HNPxEn4h
RYf5JzfAUQjCurlxhPYalc73G473P3B5gmowFN7wUKSdPYlkAYj2O0nHE9dgf879
VPhxtXQyhij+jMfIVBLgv23AZFhfSpXyUmDmJZ/lowRrRA+31y/upBvZW917nb77
D23vXa9KJQ0eq103PfPcEmlaJfZUcBBvVnuuPJWORIvWZgC8yp/KqTahuSbTid5i
chyBtIx98hlV3fo4Nld2gdkfsMTz/4ThQHH+4NRi0X2QwKRDGJbrHmPomWdTLpoA
uGMzUTi+a+zVOQkyUssxkYXxVqeX8Ip7Fw9VBRufQtX8ZKn9HujtYP8/Rsjct650
7BrNP8ymrrH3+2cUTbaVos/v8VblT+5DKKJu1HGIjTcUEDO66qjisdRDquWkVRhO
7gf0sCN77r7iikU0ftLkjVjaCT+DPQMP0xbwkRoRZxNUsaMu9Un/v+Xo0aHxNc8g
jCMWI2CaOPlKwaO2AbulgpcgeChesNJ97e9ExfrCThp/2551O+Vd5qWZoXCB+eKP
u/2L4eX/de0qPOz8AERJ7s/070HPD9e2t7VEU268eLzmf/yavJS4PFJChifVs34r
pr/S5su8n0vtPMgOfoB3Xa5Dn9VoI7VpGNJPKKBJPXQeV8AjEL81De6aaSxeI/BD
GOJTTN9+D3f5w1NVcdmJQWBbq6ejyR4y/PnqrSJPbaDzjk5VQ7PYYu4fSq5foqub
3IvOdIyzqJV/a+Fzo2OqWeRzZz13Mx9QcNLGgRP68kIDyjjpbTq8BW0SfXXzmr3/
tnUhT+YdV48oK/2Ws6EI8GlpZ55a3jupxn+cXySxI7IHEEQX7y98QCpK0ri/yhjE
fluCyhtjD99SKtkp7Ryrod1Yx/kXG797W3OSKORXwtU1Mk4nQp7YXjuUR9IxRXcS
HvgNTx0r1JA2Z0Cz6Wt9QbC1FX1mpjthSc2KbLPnh/p/z39r1Ke9siaUCIwlIDzr
idhXR9GP7aB6hidPkEYQSAiUyxhBmqvbRyIdkzCs0ObC/p99Lp2LbkvetMso8keQ
VpYeTzLPnPTWOB9nlHO0NjyIr7Z+vuOLEwbwwHDqvrQoRXXxnNfe7xvL391mUqeA
cFrmal1lXPV8d++cPUKeVuSm29KP9i7VffC9YNVSNPRfmm6uxCemlsHCBmlI6R1p
VfPEyP5ZZ14qnb7wo/kyzqh8Y0A/bxJmgcFrCwZct1y2ySKSQ44LSD81ijIl3Fwx
kqxC0xmCLJC0cjzvcv6aOTBEzbHuHODSKs21IbP/2isQZ1o7dNNMIXEdZ//iassX
PYU9klGrN5aMQVLr6K+MeD9ylmRGeCSDqHWj/TIjL789sp80f7j4ZWNTM406Y1JH
MBfvb3Hv8gsi4Hwc7fRXzVnaSmktk+gxynbHnylQ+oUEeE/T/ykVSatgM4M110nI
u9tLV0QBb4y48RHgDF4adTQ1bq8jeDdvHqYOx33B1tAD3K4Lw5CdhI5635l2YUtB
GImPIG/YtMIz7+3ne8/1PExVssGuFTLLI9tdYiN6N7kVedjUi64uhCzOCnfQB390
V8Krq+BZXivhSDPFXnGmW+DMH0JYp695xAaFUQDSZaxev1g+ckBYwl79puKC9NO7
pzTcjZdLo2MiCOJOBrRFXKw32u4zAN0NgChZZSdWgV3oh91zOEZhkZkSDXLlOFL5
NM85WKpLS5tLluHDWNs+INLTmHWs8ZJ/1YeXzm/gZSmoH15cXny9TKIqBgMDAMcc
z62ZXHf8avY2clkMIqaxBhyC5p56fFMRVFLjafRelCL+jlyjQic4U4oMzrqeE2qF
ApJcsAN4gEEYLia1wkuH8qcr25/uIeGLgjYNdGueQnfqNKse4XVopKC7rKS8pozx
mkeEWE6Jd5mrOJYlVCHUqm6zXhJof/JY4tQ6RnPvZ1rqFRCuWf4InKf2OXSqTEJP
CpHa1nnzvMv4zPLV/0jfmR088TD7kjjkbYoJO6kaB3olQIXDX0TQUvasU1Rk8aMg
9XDok48c7O8gyAEGhiNDwaQLs2IfE9fzRLYkzYNjjjSs+YUVH/3vKlNalfyujE+D
XFPJW5GDMjNojyorzhSdUYCYpAMqZhvrMHtMYacUREyFeI41wvf2LWFjACBtUXAw
1D16zDcxH7uGqpADz945k9dtr4JQmjT27Rn6I0mF/RuId5pOiXSrKZFE2eskOu75
tPzLWIM4LxQ9F7Wdv8Jyb2iOjC4HjCvPpaNRnOnC09XC8zljYgCC0mrWOEBy30s/
Yc3EHR5r/69BtWNkeWtWAokjRxAV+ZgZWdpMdDVj/viuxSQPyqSZg+cTEcE8FPNw
JIPQkqcrQn4cqBUOGzybZHy0r2QL01/R/C1pmn7GnYyDCoyPTVKjiVCnbiIGaaHV
4pqdpehy3S9559XOuuYbfhSzOtFMZTNesdSeqqY/JhExMTWdl7uUbYiVEZeYqqpB
65SUOJOu5H2ncDJjJi7dHw0/mPfs0H4XRe0+zYmBl4hLX0IxLvtiX3T17Q7Ktoie
+P7NaQu3BO7kHbr+Bqq29szOxLfrFy+vVjHkVgB/+TOuAlBKNrUmV1kp29km9Vp3
sowNhbMtX75YrOU3GPpVAiLnLq4pjdbYM+vOA9bZvrJ2Af+qPNvrOImvRlaoDmb+
2OokIaNqsmO/KUFQ4DxK9ypAFSa78Xony5gJX1xZJFpb7XlzKNvpMoM+eS/TaG9u
Wgex1YiCWIX8XBd9FBZm4MQvV7K6U3RFG3VMLL8dkmwBEl/GRHGd3NqSQh/NV5iz
TidVFk2a37fmMDZJdNa2vdf1JK6l7MC2tg7a5jm8KOYUXG/W4luXq0D7MlcttrER
K9fWFuOui3HfGRR63qAUhFdQ19uP3taY6oHpwgKAV6hnDVw2Pcg3j2MApPOhH0A9
C9+Bwo87V4v5Wh6eDGVytIqitSddlEt61zb8WcYVyHZVr4s6ZQ0lGY1DB6TnHFA2
gHnFJDselRK9RLM4inowMLHsjbho7bCrQzyqGWpwvQWMpg0nIOtu/V2JXpSOVzNb
GIMx1lE3FIQM928hp//TTxYGpHgJ84QrmO4gZhEN8KXkuzE5x1i6x6E6NLFuKHia
wM4sbExT416Q9NjWQSb5gY2eOdne5c6isYwlYZZx6sHGWfJ+Gr/TiT18yl7iFQxl
1FL2ei1UFJltNvDfcCEUpf91tgTgHyeJLLw6sd38X83epwS2MLM/eNY1onVWTeIi
xmjoPCQKY/GyN9eJXnYeJglxpNvKuzEDV56lcRLuBpS/V6KXQqNaeQ1qX5sNWPBt
oE1DYg7ROj4xATRSxMPbdTss9cUGmRtcTQt8UsQRKFsSohvzvltUYgr0W6Yqvs1Q
7QsrZJw0zoR10EDNdaflZqdrZj7hCEW4cSoSARkN0n1743qRpew70I2iR7yo8RB4
GHz+WLx3bBE1BTkEtWPTnx+FuNd6sxAphmVtnoAAsGa1EcCXXo6iczjKQaKrG8Xx
j2ZWrN8R5Cbjv78RpoLHbxpzqKkT5yImWheU0Bq8FzGirYIRpwP/VY88KdKJY1ns
AErmbKHVAF4jtHYZkCiMotEAU5zt/QZ6jJMbexr+CbVQ8HSXZZzBaLWm6vi8XfHE
7WboO0JfCRml3P3FTUbCrxXl2IjirECmnzoN+OxzHBlNgCfi2bIDf4zYarce4A2x
KBPRvQ26/dlj4uTAwZGB/QqcweaiAgrsN1NjbbWacVSOQAmdyVWG/w+/bsSnAqNo
d9YK2nbsKwDPlXqMXqF3bV0p4nMxvwDUUDmY40bDCAYkzaw8r1b05dj5yLnVAeIe
CsAV5IPFMylR8V1TjHQTZY397wlvbMCRkd8WN6PI9ulZtY5lX2sOs/dtWgp8uhQp
YIjcGXhXMLqyVRU2gr2ySRsz9X5foDi5Ttf8fo2pFVD6GKsXQWSRMObYalFNDMvp
njF/9UKZnUY/iKlsPbeBopWJZ6TcTTcmUNyO/reUjaKoU38HwRrcYOp7zArBS56q
sCi6C/Io4UPznC3h1CrF2orsNyYjZqE/7Tm9ICIlE0Rut6p3MCNJwHOF1aMceKNA
g6H+SQUOFQrPXWS7aCyrbKyJCvjziXqXG7Z1tHqE/oikimmWTgiA8D0v3Fjg9gBB
idxGpYQkqvVjEN/2NjjNOa4vznSos8dfgOzvUpeyqiY377C5RZ8dnMyZDBgF4HK8
FIUVc6IXHF+A+OfEA9EfOahAT1e9zatv/imdYEAyUBo8snJ0r2iTY3jecRTqQC3K
mRcMXc8UBg59Qc7MbilE5PJdL/6clBJONjruELbWXfqKnhhS3X156XWQAWop95Vu
2NV23sRo+BZ5QhdHznkVbRBbAhc38yR2iQ1UlJ8wBBemHH34KdihYaojeVX1CU1y
evs7gwYboXIqs35FgjmPdoMxmlV2Zt7DbwPB4BK5iGhjziT5TnlLHzT372BX4apS
OIsmPS+VUdigqX7hiiuJK/spa7+XSXgMZV2V03wVl+rfk2zE8ciiLWik4+P1Z5kj
vptJOg8wlfwnGKBxVeTXk5xdZQwYo4pcjviMI4wtrR7vtnPebh+VQc1PcSrWatMO
RTCecyxKCGO8wCH6cCpT3jEZoHv0T/U04phOtaMahWrNg28Tl/VUfdmqaQ1wP2W4
Mli9ViIlEcpIJ8jdZ37yQYBABNqgJszYSR0p8remHCzp8mDEN37v8ZFimkzqm3RI
uWJJmvDklCuJuGcHcQ7Hk4L43ILcK6TTASAeiku2auAGDNEIGvA4WKQjE5UhYDdS
N37CvjES/IdmVsfS8m15RKKhfzbfpN8MCYdb5MvAAbqwuy05V++26bzHsLLYl9ME
v38VPaD+sK54LUbQ0ul2Kxxvjj6nKoB0KtkycwChH41cEyxZ9+E1VR9+28ATkwrm
P2u1MtGPuJLRUJn0DBB0GLUC6vShuqUqTomFNPOOgG8TvH8QwDvVxIPcMuk299vB
xu+0uZSiUBgz43cqSiO6UIO/inB/no9ZU1kieS77cRnUzqj+kgpVGP0TKENIYGf1
x3tWwaYT6M61+tiK2oaZe7Z9RyfkAF0tW9xxl2NZe8OXaYQg1Ai41grTVHDQGgCD
JTPA8umM31iUFqn+YoeBQ2vOqaFF6ZVRox9D+jGXSf3WGMssWHCPGplkwO+V0m5X
XmGhAFN9SZt6mwgL/g4vgmQ8in/sJiDLGIaf7qJJWA2wsaoyjv7dtKyS1AL139Kv
jgk2Vnlq4zndn538Iyy1SP3EL6L9GDH3X3xn46tqGRQnZLCRYckdnYEAZe0u4QlW
LuyEWdWklQ8pDvdep3EPQzD4bWICAg2Y8nWR7LFz8BlGS+bKdcN7oO7z9TOnduKC
31pMLZwr/K4u+kjwYFdsBSjey9WbohBjGCsRLZgOFNeFEx6uzYLvRAw8Q4X5g8hQ
2b+P/FTKYRkXtcT6JxceJZ8VtzI83mGADOJ/E0bSUExzz4TdwMD5qsDxZSobZyHP
jBTlxFAHCV88+bWG0N/psxAPD7Kg9MbUnqC+3/YCRK6Yndwmh8DAWyIJaooDbpu3
zCqHZ8ib7xvqZnUfyIGER1PLxpjKMKM6iTasGgkehj8lAOhQMIwOA1DcAW5XDsXs
juGeBOGVFPCRUQNa0CUwd9gXCWxBPltXcU5kS3MRPpBai7mZ8OXKX8Ph6Djyf0LK
FCqFo1PIgxYuBHo8ZNerSzlldrRRDu6sdT2v1s69Sn5wVJ/qMZoACMi2ddxpckmB
gtygaLJ8F1VKKat6D/QTILC86FCdM3UvTE9ata/SmlerGFSyjqKIIjmiII4Jx7Sz
rVeOnGbi7LYVVksPv/KmCZFmn5pjPXypNb06e0x6rn8NHUJgEF1jfwxVd3DywfpO
rfoLxI4X8HcV7SG83eFNZvFloRaBeUjOOZkzqvkbCe24sqEXsnJumPAiq478Bgyq
StGpygFfFTfDtTx+cRO8js+ov2+1OzY3AzAG3tGBXRh2LaT7iZWPWqBagA4nvULu
wXBwnpKmDm8taRfHAm6SdNbq/G4utmrIxTqddIDrnoyBpKKWev3dq8J9NscJjt9C
CnLTYALv0hldmY8HGXV8pwbKFwiqeBXHmwHcDWv5jQgWqN+lvAq442i7uo0qnPdg
KwvOpGuCQalDJa7OrVUcO5TrfRnc4uvtxhJym/EW64QXdtB/8r1vVNDVZ3snqH4P
8iBnggJ/xmemD9lz+/6lv/8P6uRl8reUakPaM0tWQHY/9z8ziwfybjcvQkrfoIuE
nKQIJ52Q2wIUSsPm+8lHfoAyh8rM5tpLjEsOjhrAh7X4T3BEs2EB74sLi72hhmPE
rFBOoqFKaDS1UKveeOLY/Von2/oPfc4wIJ+DRA87ERroN7lyXFlxdz4w7VaZC1JP
GjOvK+F8a0IyX4ISF3iBwigBZL2o96fXIHIN6kJwINA1u2OmUGY45mQmkpQMQ2Gj
roedit7j6/zWEVIQKD+5c9qif9DaX0s2+xnJ/enFIXoab4pFyZGu/mW9S+15/doT
RoGUNETloix+irbEggxOfvxQwER2YD9k44rERMtx4SRvycCSmFrTSBjlyOAzrEaP
Yivu/filQPV4RocJzzuAfeA5qL8JA+O4QbqfkDBVJNRPBymAI3NnSxrVOZSwRk7o
DsoS0G/8lOx8cWyYyPYXbWbUvATKHebRcXmWjJb0DJvHnwBS3Dq67XggRbeeUjGe
F2Igl6CjYYv9eFESw+FV8lrLs25kc7mj++YKNPn0hQ5dllPhX4+l7FL5H5fpR+6Y
W0QHlY4tFYY/+RHLF6iinU81DLvAve68o144zCcINQIAgclorZRemDCoguj6UlyA
QPjZe25V+AZiNoRURfdpnhlH2Ugr9L2A0HD9VrLhRx5cpSPz+X7Tuwh9iwXz09bD
u5MJv7eLfZJDJLlrrMSvGkR9bEaDRl1bzWNuYJYJBdwbB4J+6vY/+5QIyiRkqo2f
3mf4xD/V85gZK+FRV5VhX2YAnYTvfStuKDCL+D8DYIn8mG92/rDPSGFRDiXG8A8/
zJEWy9yxqPQHXZaN0VXumDOtJ/ORQbTIqcxVEjGC+Q48ZuFrJ13tcqAnUEIt+1RV
O+GFJg1vx1Ne+dJlbHiA6Gc5MDL8I0IOQ7dMg1oMOo7iStPiZ3LcfgyisdXkYoiS
iB5d7eulqM1b91434z0xJD1z0i4H1U6/+DPvyu4VAR5199Fa9ywQb6UWXgdzlYgo
PiF7y/TVjTpOsuElWMvhIWS2YMjpini75UxHtLEosydMHVF72GShV/yeQ02ZZuhY
2pZ34bwz0BzSR/Lntqi8rw+5pqJduwnAgB9xcexbdEJ5r0qJO9jcE3jAG6dSucnJ
/CxtPZKnBqqQmskfpKM1ELmwy1lVhVZczk15WeBemZo7O8DRdeAwUmELpardT26q
FL8rjnvc+64C19/8saU/74zTc7zFAqzrgO4F7tA0dph7EnHGbvnLJvah97LGWrGn
xzgi3S00ifqy0EnPuJi/sN6zTuTA+s/I9pCifxky6IcKm+Uw/c2wTeo0y0iAg+UR
WQdc4I2qxgNxibKnuR7g5yJVWStYFyG20VlE5E85XiCJdj1g2NuA+n2joStH0fh2
WH/lkeg+ckwlRYu6ijBcFdkugSirtcoqNGaIEgs0YPrtMRZqA4XutmEtRepBWgzD
SPVbZjy/eIG9kUMsYjkcUWMCTftRZg2ssii6ySfIXQ1sFpPxyqgcaAVwL2hTj/XW
LPm0LiX+PAAFkoUv2Tx2E0jQVwjotbzu4wWimiY4VE1F4dC6nzD7trj5D8NIyQ7m
1PHOQ+MBFqyuxVbown+bbqdDLnrfv8j0b1liEnhA6EhbPUzG7Px6PmuCTczavLOE
cgZmZPW2A5TjHIB0H5KLzg7H5oDUOpAE8xfURR0si3qFRbrrU/4iIgSwxB1ZoIx1
LyM91SKLu5DhJEv85bWHKMSpC0RasVyp/KDwGO0vAk6wzgs3xuw7i+1CvgxerQZQ
doACIcf99E9N/GMDRJDFbt71mEADcIqDAzPXG/uGz04PD/fsC2uGkuMtPk8/9PxU
DMxfp+hCahvr3QlZzqa+e7B4ci76p1rEtWlmUe7AwJQXD646R2PuHg7MoO0psZJ/
xnMXAtnsepTdMvIDXVjeds8H+tBcVyB0d1rQqrOhbAHUaSm6zN6F+92TWuUUhowF
rs9DQuZ30+4T41rS7z60YvGqSeeaNsRd21eBt2S7AQ0aDcwXWV8d/j9rLXf4tL2/
Twh58pAbq8tJhtR9pnwc2lIY4ecwtT2Upt8mNsThQ7u09n5vsczpghIp3UlLt7nN
PRUHzekNhYMm3f0RaRiY8jnyJlC2rbDgSLhb9WW2dKLzMnZ9NpXUdYyZ833Guong
duDgQ0g138AFZtgXMuoji08BMZ6LsaU7Ce9bsGjcjrYfyT+HXgdva1n4X3SO6TUN
JqLhn2ReDa1IUUm+BtwkQwhaDFkMtlOc42JvUQhE9IvXXZgQztiKiZBmAvagvRJo
ZjOL9ub/n7dtekKvPDKfmH+i/JujxVjfVcerrztuKgz1n6Qn2uN4CdVptyeddMXx
wgeqSU702+Dp9NL7luTiIUH24t4cpmAtG0AMs7ayw6xTLSh/PCUb0bqACM29fQxP
zYtbz/D4PKnuoI8ZxJTA+hSwEObxaLMn8/F82KuEJ9IBdBFsV7Q52GJx8BI3qplI
39xtqmbIVe2veGs/QKSP85+SJTk77tPqCCsGepqewJagQ37tr7Hb8emhJ2LdESNW
RJiZ+ve+mOxSGY1GHQ43xCJoWvHVm2s98uP8RherEcIwiqRBa0rzAj5fF7+KIHB2
O28/9m3/bA2OiLjeYbyWS0bvYfKbYbuwXm9iRC1HvWwKdV9ZwSdNYVJUKOHTnd6O
Oepbl0l1pwDXTtbazhF0jXnmoPhnrQQeQL1mxND9y9rXdh92gG65ub/IRm9iuZaG
2hJfT4rYvLv3+VmNK1Slbwz5dq1nJr9s0DpcVeQL2f7ES/YUaWUIQkKy5TldZXo4
z2kQoqd7L2u27KqBXlZuP6O/Hwg+Gf4+ml2cxlqOTQkSclQhG7BJcA2jZuEzBdK6
AJFEUPIAD7Ex/CXDtdKW8T8EhRi3t0TL/QdR+VqryHzzrWIOzqbvpl+YK566LzNB
dXZeQtactni7ydN4b3G0br18y/EPlPuZ+fiUv7l++z4QO9t8Z8D+ktIK98rw+VC9
nhdSwe4e/SnTg4V0DK6sKQ4pv1MnDIlzBZRPC7HxI6Fnq1Wv8Z6SuKKskXI38yB0
h+DbxvRx579SgRNC5KnVaYtdkbsyRNrvD9ijfMe00KBrJ/VHhbPrfKlhJ9GgIsEB
y1KE6esI+a/iN5S4Zm3LVKJAhm5nzoVa+l/sSzNA1P3fwP/55nnQr9eI+LBoWFQr
A5cr+7ZMq5tTi61mMcunVI6xhHzw/6cWI4ZKUGCPz12mF6+EZ9tNqEMoa399mY/M
lcr92YCTeCtWb/xEwmWr4j4QhQh/m/WSpffeTYobWICO/U2P6RogKSEHK0e41ii4
X5qBQnodqni7eIS2C5GALeItvq/N2Brlm0dU89PTCqfqTA6XBTJBf12U7+p4U2+8
7tX1cUUiVN2hHOe+0a/FB52hQ2lLIioJmyTpiJ6C/PMTHyV5PTiyl819MrYIK5BH
cGK3t/iXswUkgwBKNgz2TsVxCq8sHMT2ZZsohhUiYXPCJjTozraD2RaaIOwwFNM7
eSOYKxUJdWRRn26iGLtS25hbIOv4pJ49mNhgQ0hdMbmFqQaQFgBN7LfAOb0WCxYE
4KXAr2QxirKUhIJ43ZfrIpcVHC9cuu50JRnT9oa/TjqQHD1KAe6LeNm2xj2aoH4A
tao1uQ8ekRWU/BZuAGyRHcSMRPE3a/FSz11PYdV9QJjMkRA51yUT45yZ4i5eDOZp
zxIKmTboxVODHRl2akYMCxppIZXK2hX3SETy0P2m5EgLsPyX+osziFF6/ILFiLyM
Ok/WX47Ec1unNuHtyBnBFmLwnWel9JFh7NqtQ0x1xr1rxgbWnrJbjoYlhdWcl5vy
ojb9qM2hTtqGMiRrIfvXVLvGrGr4yjb5VkvnriKn65Mkxs9oEvDgsd3VBmO4zAax
X5n8C4V4dN9zZjoDnnFxRzhgYraiwVW44hB1j4KPqZZzNrg84fHCPVZ02M3Jk4n3
DI3JL+TnpGv8e4jNZRWJtyc/KOTmPMxJNZDfcWxnv+Cu9RGlKvyz5NIlxkCNmXqp
iUVvDhA60hTrME8aoiAy2q5/bBETq0xBzsPHtt6cF6TOFI5vkvqrOyvieWv3ER+v
ikAMz9mRwYLY6OrmhFhF+MXfkCNHbSbOFBbB5QQB9iBYkahBx1jdjXjmP4blOw1t
ESsfH3CthUejMDhQ8xXKhfQozGyoBa71zdlt/qYxk2qmaM5jwKCsh3inCOtr/CxE
MXF30Qd77ZLXnpiSuQ5JaSGYSZYkLVAbXOAkYGMipL6RxxV+UFow4GUTuB9m+Yvr
q/FM5q6Fy0uAhgyr9SVEc5XC5Kv/a7pK9ICGdo748hUAAscoi32Gvhoe/tusDFXX
b+vwQZqFUsfAi9oieagKb5QnnduvnN/lHcaCWVARAKL9SHSmfvWz1Q/W+crHzkZo
xt9PMQ1U0lRlcN2Iidf6FyCZVJPLCMawz5djd1bDCT7Lep8FKV7kiWy/e3B9WhIr
VtxTC/Z5g7C5+9okVw01lZiHFfqJVW3UwuAsDjaiYrgWMfmTvq6wuT0BxeXTE95z
KO1bEkHWEGOWXYDtxzW5wDS4uppGB9DbSGLsXq49l1DxnmFEZkU+pXZPT3pB/Mn3
BJ2QJpJXy0+ME7zYfKQEjgU5oDdaufy7srpHLIkbhUcZeF3WKoHRkrHr+Do0prWa
DCtn5MZB2BEq/tal/NuN5Ekq4R5ZDeS70TF1vSAsa1+LDT5WYzuVkmZESWhlA7rv
fnqYd0yVjI0Za6p4135AxH7TUaibuD0Vun/KDRPpwxuGfwHj3cA2ljJge8piCi7g
QziPLSLl6Sfg9i2/6KGP/1kp6oTqXrINmpb0/Q+9NfCgmf04prFpt3FCTmwk0vlI
J8uLhiad+edTwzXBt58Co8kjP4Yh3E+JOTJi1KiVwv4cH4zPkjvOJy+dI2r6byYx
Fr6IbmFkGIkrzMxv/SzQ5CAl2CElWNlHEVGkbakTQKSzoTNIIjfiUdcl18UTUTyr
glORuc4VoszWJlQ3ezNCJlCHsK/xdKJjb6Mb0EabyQlDRDMQ5PtIbp3lmr5jTZEj
G0tVds65bQs4Gxof/JKh7kLWDFFdcp/dPUBH93vlWb6/+6l7zBx2AzQI+kUMwt8A
g23eK24eSOrPtls9QTH0iQX/J70srba9f9/Eu7ISb/lNQWO3eKjX/pbA4u5zBwjy
Yzc0Pg6ZL3knM7UuDihcKYCvguhWodW/mhcvHYyq4tWRIDIcyTXEUZghsjqfzOmL
YYG0uCbF0leksXa8W0ifzVTlFJj2CCJlqkLciTTOnDoBfP5dZUCWppd0mcSnNoXy
C4dXIh7AZx1rnDqFvot/qHdjj4392HHxHNkxAlfKQ9O5eB5By9MfCOqsb/t/yM6b
HtTf8ZhaO46fPF9dsOno5zJ1e3TnOfy0KhhSAbjebYNsAUG6sxNoXN6TtmNCwbhf
VEFlxq2jvuDije/xYV2qtaAXA0Wb7mvdQ9Nrcz/LPj50KRXjOxG9gLQgTV9Cewcv
Kv3hFEl5Vq5LVPhcDasf1XWjbGJehFO1RrwAqbiC+WTYsAhr1m1IkJRf0x+Kb8Y8
vSOGo+81WS/UJVA0A/g/OOP6N3EwUbk7Y4UWS1dtmpl1t0vc9j8Jc75+EjYXvKEv
XZ0ylE+XMsV6bDvWDCTSDNC/Dk0TQwUR4UfETJv8wKF7CY2bQCLyGhs7m7k1rw7U
7RAGBnKGa9ic8b9SzeM5CudGKyaMf/WLHPXWZ2BocPArAw/mPr0LoM9/jMbz6fzp
BVpqu1ZrmPGY9Zl+LaSNn/c2284Q1Rzh8MhtU5fEAsospj2VtlUyAWUykxr4WALs
bEdrkUoB7hHxBG3NqvQmffnsMeXfAKxntU9bhOGXKKhXK1MVTUGDXmqVXvrgeLuF
9xOCsOqqUq6vkoxSdbjfjRUQY6Clzi5x4QVl8fV/xmEAI1UuvWw/2NMcDoGrUbFP
/HH/QzMhWvYwdRveZkQugCHJra8VudJOvp7t5OKnhVBlVE+HlPApNcETGKWabUHF
Tyw3U15cHw939uJFVqcbE7nS1sHJD4ErxXdsPqreWUwQteFWSLLxMceQA2+TR29B
OFe287DhJ6YHXSpxhfsa5eNgIIEHdhgltLQzWux2oPpQTokhKDXO5jVgC71N9np6
k6DcWXFRWA2ZdHAsxTDFSNFmC0IjZJyKS/mm5y864Jc6DnkajB5JhHCo1iplTlbD
NjzFbTf5z2nrsONCQZZkTQUNUk4LvDE8LZsjItPMTNRvLX8MfGe2BoZLWrHPfXFr
U2cbHCjNOfVUIq2CQCqSvToauySVTJz0gSqfEkm0YOKN2p0FSY3Go/CF7TZRvh10
3c3IOzLuQRUjWRVk337ouEoOkQNL/zvEk/P7u8l2zrV47MQ9LwJ0qsnnrFYTh1Mj
WF2sYWnjUw+aK8LVB20WewTRv8PjkcxspXfgkyIvdwlzivj2bkMK76bJU5pYFyYV
3pf0Mf2UweyOZPB+OwGtNt5y0aioFYJVeZoIgUxIZ+3MVXGkHovUEowONvkhZ+3P
n/syJZ0+KH4Y4Z4g3gq2RGVHQb3tFKK+DBp4JqU9P8JgwRlyq2gn5BUmZmkA1W7I
6SRfvMZaY+Ygs95Ioxs9HuYMRy/cb6SHqsjKFrR5q46YMF0pgFvWkW3ASF9vHahl
GXWMudqlF+zmAYfN/3oIQHKw84e8KxlWb+sTy11uOX9tgHGdSxQRns9R7O3soIso
1y2No/1XI0lbhpTMaODsdzOGZVyy4GrnUVMTWuG518jJVKX8I59Prce1UorwUj/W
j5RjKppBEJqiBTnl8v3miIsuJrzWluNpWkWgfA2tLU25L4LHYr9vsXo0cF/YNzJ8
085WVaya8hbRemy3+wVphfXaA4qWJYz/EGlP+nzjki/053DKPGUuSDhjm8lJG2Xs
gE4yOaBX31YS5Fb/4ZA6ERLgNkPcCvqJADcscjoeD+sSQWtAWe/pgixgoQT1MLJ9
+DWlNBku/WWUb2fOnFDVZzOT1cuGUTSjfxOhdg/phcw/sk6kT6FWl8icitYdj3rC
DTVL7TyMGhBO7RwcykhiDoWi/Ok9wdKld4NRguBlew2wVT3NtvThGBJOauW4cNk8
Km9eT3we65Ur+Z5CQFuY4J5Ui093jxqp4ycca9zN6eZUO8uFVqp1Qvub87nfv6YB
aLmeaTFLMG4z+xGcrWrIw+R0SC0tImzoTIvglz8juo2AEPHHnuweQuMCARoqMMe1
L1VnseS91V41xb2ra+G9ja33Pe6yOKykrGLpxPXHgw0ybcrhjqKBFL7I2lWK/Vsa
BPvYjwcSWtaN1AJCvfEotDU8dz+Br+mHaIRbH+nT9MvgYBnt21vbPgQmFs5E5sz7
PeU/+1ioSE+ZVLGoWpD2EMDgAdB2xA+LUosRxjQyrfeId6U/XD1Xlpg5lbwpV/pH
+s/MznV/ZC9AjqEMPZYZk71ccnO9h+bIasAWybrZwYlVvd3xBu1EZB3zoK4KBNVQ
oGiGUQDDH4eyvJO3eH/Vzq+22wbLdZBnLgEkenzqU4WpkjO0IGisMdzEDFWG6VpM
SoNmbhSR0TtPLdffnPls0WFlJYSET59MNt/zW2+nGpaS3EqGurcOjPB4AvnCS/Da
yFSw8blyjw4Zm450FNig38SgfnG6HB3avnOkKiqsE70nC5phBQPCKZF2SVJWTZ0A
Cx6aICq8p2SIlxI4HoSMV3i1U/rIjD81+bRSj45gbIRACzT9+TkKx2AKogbpbDAl
OTc7UlNi94w1NbBlyaNtZxMqqFHO4xc3+9d0ePwFRUmfIB4kWNiBJlklSHKE9K3P
/VI6pJF3YHkKYRBIG7IUMEz9HNP0SAKeV0EY0Pq96cE9DaA7YUvE3eOLNU4R4plo
/UPeVSDpxjpWQnzDek5axbLjctVLU3iMrXmO1AKl/aacoqtl/eRncSlQSt6rxEtM
FbJb7tKeRNEEo3eOrqIB7en5LSbmyp7qCQOA4vEadrurtoRFO0JzIV5BfXamqsHA
D9tl9+lQjqchzRA1iLRvGFhb8BnHvIarcrH2avYZu9LwinB4IDoecS34x54WDNlt
+MJN4JjCfZkqU1PuDk/QQJqxajlMJwSvKOQ0yKGFwbDByOglm41lLhGwwIBfP20s
Ig8CkVnOX4mSHrNk8MfolTOXgWOUzQH+7StcA/EKMJAp61Ko8GJ0bDqviVbHriIa
GKjcMcH0I/PuG5ZBg1XQcX2Tjn0nCWfopV2BUsO2GjgOaS//pkxFPX/nm3OaVGXQ
os7TP6PyX6yAwYMxQxih7oqg0axEvRzs3t+hkSMtC0W5Wuqm05pf/NFSSM8Za1qn
ms0SAnVMc7PS1498r0o3AhIwQhM7KZcZIX72Chvk90qg6PM9Ticvp/0K8DoSAjr3
zmIwW/wIzY3rUATYSEu/ZVmAY6TXLndLxlPE1ghSnSu1KtPHtzN44GEhqfKgwlqh
Y3sQ/nV6KeIip3fwWqe+wZPzmKBaFe8nV0D7sc3WJ54qCLG6tTC4JmtatoYo9d9f
yeqNchl4NuNeEnbVLxP82l5NXQlTwq4WBOjNVlnOXCmkh2tAL/V2eIRpTvk4sLRu
6gmcbng199C3gZ9OUP8rM5vWPiRa5yKAN4GQ6WVYfEYqP46IvMTaARqeEbBnxw19
I2Kq40+dtYmbXyXjHQvZY9mQmXvWq9/gW4p3JrYHgSwE8XopjQMfvttj/CUq47KW
qX3pgFLLRocQeOkf5Xv3iLpFzy1PgPrnQSSlfGMdpV4vYpJDy388yE3ekOqyt991
kQOwIPhZ2mALKrGAIrond1/29xTKdm1lvWR7oa2gDjcNKrNS4orxhmAGn7fsj75T
9kssYdnMXmCUVyPKIb07L1ZzWMi1cgP83IyMbysICqw5Pdv3LZRDO4jLvg1Fw9A9
CP8Y57Smc5fQCoFHIOP8Pd2xyX7uOKId+S8HrJtwPyRMITUeWTcB3+fETUb9LDsU
N7G5dTTXLqOayuDOOq2hmKISP8xLxJN8/1Ok//oViiRKM/DXaye4Nxqq8hsZNdbM
WYLW5bAjzEZsqXJEHPj6Tgip5eBhXbRJ1omxlMlSadl/Jw+y1QFtn47UzyMOozrF
D8qRQLeq7LgDF3ioz9OqznPt6GKV1YaSJAOfqd1snbiGmwaZpPTT1KM252CH2Sxk
okWyY/l6B7rMRNDsPmfgmFYM3Q09xQGKl+OMtf87+YWzlGgkFiOXN8dXDBZ6ohvQ
w4eYJsD1XBtyDWugiYKZ5X0kTj3s032MsGr3VMVlg28Oqfob3NYA7bw26DMPMoGn
uqyc5hK6KB1UJoNYanbxXsuMYjryp7bRwZxG9YwAIuI/1olq67o+JmpuZ4O0OFMv
H/BztwWYjkuQifnpnd9yJvE+QKocH7QC/ftsFF6yCnJ5B+Hd/xBzyJ1iTfWvgFmB
bY0PDhzlL7DQWAOl8LppSxyiR/YDlQbXwsN4T3p6EPtuxQ1eerXx/vhwAPmx/NDx
mFtXVDG3bhOj1DDMqkM+Xy8AfqZPIrln0zM9K98NjIzyDVMNSHYDoHq35SOHmNhr
6/GWwMk9yU44egVIrOwCWO1wzS5vpK2s7oqFydtJSOhBpxqcA42mJVu/h7BxEfrd
EgU3acIIInacJb5vPLMnogt05MQQjXpFr0tvQifW9PTPg+WGVDpKtzbG56bB5VQT
tHniBZ8ry3qv7g+TAdlD0thJuzcyldQhtm17eNUPbfs4jNqP+VFPg/HecduPtBZB
rSNyxYk+h1RnqcgBmGdPEOPKVzFbuUC4F0O/MMUw5Lt0nXk9/j1PLcw6i3yyh5GX
xtSRZHcAD68Q3n3tK94HcdGfdpt03UMNblUfpkvSMacmx6mRtrXUcECsn3GyeXhO
koO3vG++ABQhwdiw0/7wRhqEyQF0iOhzpZA/NqAy/XmCzgjea86xo5nyg/ogxjHQ
r7q5bVQMDWfHs5d0ydvZVqpkHuFLe6rGA8Q3n09u8GKnXFdM6LjwzI+q3c/Q9lAA
rmr3xoOWkQhiH1xfq5z3cejHHpVRnWOJyJdYLHK6PWqPEx9PugZaGiO3Dr7bMUQ3
LTxsTh8yFsPMHCVXXvx9aaJJe5behX+MACask2Vb29oVo5tYbSP8T35W+AdsGFhI
p2MoySCWbqABOH4yHwDGSuhHZsy4OHrCQa+H4t4sprXRVBQsApnZXkxtx6Ar7ewm
I8g5oNYtnrW6zbn05GMoubHinX6F7sqkUOSgFYEt8DMexj4/KUvgMQG18JpkVfVq
fALX8iXnvfExi3t7uSvoVYpE9HVaHUpu3iM5ORh0V6rrmXv/Cus332Fw7iePk0Bv
QsbiUdAMtO47TJuXLYnyhJtCET0qekuxLslvq5e+7cYYdDZZicLlNOSm8dfh7qIT
7Guuh88gjzsIdHL2SpPXPpT+0Z5SYt4h/AnfMPoNYIb473OrO+zsEt9JgyNfl/0X
PLSftp2yTeMhBOs/LKsfUAyvr3wZkqIC0CzO1G5RNDBCU9FPDsaisdblUCYDIKyJ
OXH3fNJI4o17xap3xuXjNoIzCsnUWu3MSdPmoJ/JwpnBZ8PInED9Ff48A+9nLUtW
62xLY+nI+6xEyhWvgw7vICY9q9SCJRpIovim71L+1E4dyhvTO3p42QHJR5uKSVat
d7x99xn5iheVVCm8cLvgTHumtD9kjuzyqXpghENUq8wswKbOL8W/gmtREoPOHYY1
Q1h6bBhH3cUCduHHHsn0VeexODh0mEOrP/b9cB6IRFcTFbitFBl7m9OzhGUsfXmw
G4v7WUFTQabAobHSjUco7Zk09Su3hjkj/1fUaytDyjIwoZ9zpdbIdJhyGRP98k3y
u5oxl8+7gziZwofEH4+oVp6d37kXe2RK1h3DiS6zykdVHiz3FL36vMfyUYvXVXDR
AgiEdHytp1m70ZX8Ftlj5FVFmoeMFSI+a4P2PieNukMazCTPiZ358O+5KkUDEs/9
jgzhSjrVBuKhLhNN+pbIJTYM/VoQ6ScpgqXbMMY2gZYPN0hjUXxWGPRmABf3+HgO
9R+V7wwlsiVbW5/MZxQ53AYdEDhqfIj+QNYzANzN8aUfSOKa1k5Nmb1gd+AHnbcp
ZBGvnpb019fSacZKaW34BgOEPDn68oKwyKk4FQ0i2t7PzKPWbRK8J/jVox6VhmpD
yJatzrY9hEVVwanG2/w6ggzpSk5oygy9iQN1z1JQmF7WGXVXNOuc+8/u4WpaXfvn
zpmmNvt9rjRwtADOyrZfjQ/wmcGwsFhid7GVqA2+MZdirZ1tA8dHjL3VYYVfVw5e
zVH8kLbdmfiwPVXuVg2cc8f3Xg6Qc1QRRtlnLXZDHW8SdwKLHPxyqb7hVV1x3RWC
QxOIrjhEDbAlZSjCrmPheYrcFD/R97h3rkbtWhiQQ09W2uurk93J6204XuhIeUVj
lh+cG3zunVPNjNz0p+3vJkVo/zg/Foxzhe5ELBVGhy2yZZkRtcHEw2IyiuMERxAa
dfnMq8kWl2Fd/+yxvrVDZ1W07fy4DyBjVPEVhe5k+Dur6eZSbQ/hKDsCdUGgped8
klpxOgsh76IJmWyxRfPba+KyeX2o0jyCM5J39MoJwd/wVVT5jSmDg62/B/uKBHAn
6+JBNIJ9BXhCfMtMN28K1jqyYE21P6W4HYXFueG1m8BSxLa2hNpl4WbMeJG9/0Pm
u1+BryAtM86gx1BwsiSsUXHdSb6V2eP6ItDr0dJvrSXrTv2+wV37I4F9GCLj0v9K
0T/QSy7B67UM1sEuqqjrhJnr+6l30T4VQKte0dXUcOgrns1rXcLL8JydLCBirf5C
9V2NnRZUv/VfPZkYf3lQTqc4FyJxErRvbLBlyA2cUHyjKRXQW/DLwauGuJ4HGeqz
XmzEv08a9VGqc6j+WFTbmdOM6TUNoZyVSGNfIXlKJB1A63KpEWWXtWlbcRh9j1xn
N7izOA7OWGHO2FqOmTEXMNhyZgopXh1Q/UCrVXYQOTKfYwMmuSVQ34Reb8Li+hcs
R0FMNgOppUALRDRUP43E98hxaJ3XyIMqktJkS6PfS5tQEPteMAxrnprHkzDEm/0P
ypAEIzpvi1B0ttPklWVJVULBsETXXespjFVvDb9fhccDJoqemjcf7zy4wgUPnmfo
tdiHdskUzwW7U+5ZT4rqTXmbEojvyE9yNLvdXMCA4hBkfFrQzcod5JaCDROYL2U3
mAT8JgpWhs1joWyxFDW2iYlJiRyBr01wUtYTwa1IEk9ZiS12WbvAsbmOBBa2gj8g
A2I15bJRkse2yw82WdNE1fj1uIltPCHPhUo5+k8mhAgjsQ/tOo+Rqpq3vdcEBsTd
/fcXnKLQkScMcZ+zb3CIZMKrgkvaHET6teWXF5xzkSZVcnLNTGVe94scFOO+CvXA
ovOPoljFGyq/NjQWC+KAD4zz17IhTpZAd5iksxV4VXtz7H/wo3S4Z206e/K35Ft9
HUY5PdcIB0oohtwV5OmSxNOYQEaqvxqnNleo+Kvnf9wP4kVH0fvpYwwjYPPAamEX
5zBH1xYzSn7O2oc7pAekKcPpDGT4xQDsK2DFNBRPMxAp2TiCbDCJW849V66THvZj
2+hqQ6v7908mtZKarICnkmxTT7q0HHjz149ZxrJC2nggkTeAbnXjgJzUEbMHzInP
XOjJ8nQfwwkDNPMZnsqR4YYbiqnyUr9ErwhaQARbuZ6Me3lxx/6TUf7g8xvnm+VU
5r1xl4vyupe5OQX1QWl2wy1AwCqLlNvPm4iltCLKvKaEYSypsxG0DzwA/adPp4vB
/rFTBmwvf7rmve6lVO6RZw2rz4ndiBtDyfs3zo3cHAbD8h93l01C80vhioNMLO9H
12hbnEndWQ8ys3TmauY1u4VZFvr3IQ8GnczqD+ytIzxVjkJyuyyU1GGfrPKrPQ+S
fummvRPjjGpbmK43rR880pR+DczJLMPzWP5sdWKZd/+hjscuLG26iB0UJdpVNBQS
NIDHpd+d9USwOTkz76qX09K9kiRnDheNTif/dzJJ/W7aFPcnFd3nM9oOt3+uoFW9
+9Q3RWyqaHJ5ybfKWh/T7FAeqIxEaJUJjpo/Mkfeib5eeJkrsxe9CHg+EcXrWjW3
cNTu+j/UrLOTHiEshz6H3IKMaVInFRcfH0UqicRhtuAiB+G7eFNVnuCSTJqy2OFE
kS2yyET1K/cQ+Ahpc7DwMditQzkmq9bX4sTxreXRzA2wv0Cst7S/8YSICm0TPyjb
QAZPBNoFlC9svsSB1+o95r8NnG3gR/rkXmvlJvqgvi275aiZYxnajZYtBR+FCnUy
hfyyJkwWpKuoINAJdcgV/F2Tlt5ccL76RzGfuaMNjk5PnOfGDiMRw3PTqaKM4Qdw
SdXP/VUEDZYC5QIktvHLmhgivo+ilvzIJ9zX51NwimEI7UeIf5tFY5E9zE3RKzfQ
Q7JD6qZcEdQBjya0piRUIIvBACmRs+pha9638CylSuiPJKwvsqGQ9+RYnbdtFzZT
0rPTj4O8ApB0ydI7bY+Wpl6IDK57xgwV9VtFKa0VSn1i2xjTFd8glms8DjsKzSIN
LOWj+KrpJSV3Hq4Z447az8+jqzU2z8kZxuLVOxBOgPLcU51dv7pEgSN6dHDXSqap
+4PxhzMKF7htOo8Rp7saaxFQA+w4w9fqYV2a+9TQuzRq0T2lpuG0lsb74WvTLn59
w8vysbA0W99PF2B0cj0QhHhxOQt9WDq8PugPMSH5ExpM5HNTAnLBIwKXzeWyOQpD
2ICyKzVdm/B7pGC4prT0ThoF9FOgnwf7FyrMCDCqVjLIatNTVxnhBEPrDUY35Ge7
KH+k0gjefvh9685u6EQFvXHERgBRcZEBUZr9YQwctmoBTf/aAjkLwx7BFOHb2y5w
CguEnkbI7GAoKyNDGb+HjLq7dUGObvK9M7u+N45dKGiGRFGh/NOOfoNFMXPccHsw
BQqZFmdMS7Ez8FMoT/1qWopF5h8172AJxGZfO4tlmkagYbZ1duyzFsmniU7pDKk2
33ohB6w9cT5qFBedB0O4bZe41m/6a4dU+oU1lwAIzZmOtlYMQkA6IG6carJlSDb8
zW8k6REH9AzhnooBi2DxFu7axUWPyDNDy1IBjrtI/YbyFFvj22lpPLDtp5TWkw2l
MLAmqy4WRLm3FEp2MardOpqyzKPxMlN3Pgz6RgsfT48HlZAK05QdTuCaeCc0ohZF
HZTlKnJ1HVfRHa0j9o3UqCyGgExow73aEA7uTtgh3T/APHqN2ZFFKhdE+HnVoWXb
twJCA/o38keCpBfUgSledJ6ij1tunmnbc5gtdDvQiiq8O+BGvE6ycrKFxJ8HazgX
uzVU+8cX3jUHkh8K9mHAGHGOzfQJm4r7ACrb46OReugLF2oGW8L03c0Zzw2YufAR
2vWdZ+O6EFd4TK2EY5LWqA5r9YeJtbTEl7Jz1HeIpcKwo1vEgjXgnJVomn4hGIb1
9XexIk7WFgmk+Ut96UwM0gQ/qLDHKcfvE4bw3b20TlgheEcwgfY6X6qb2Y49Nk2M
KqwhKixCWp8TPExf4I1BBAWrd/3s/9SXK9vJh77o4j2c7smkfKNbu3hi/Y9RmsBf
BGoX4HU5EWGv0KTtetIJvlVl0pB0Lu0j82vRiqE5hGEk79cuSqWB15rJgNekByhs
ng3qnj5E+zPs91EyP9OzoOmxLX/rm+Jk5B7AUotjNMqHig5noNgJNxi9HF0Ku7CQ
fkVBgqa0qb7uaReTei9RhQ==
`pragma protect end_protected
