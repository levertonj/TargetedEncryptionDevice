// crypto_test.v

// Generated using ACDS version 14.1 190 at 2015.03.23.23:35:06

`timescale 1 ps / 1 ps
module crypto_test (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [19:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] crypto_module_read_master_readdata;                           // mm_interconnect_0:crypto_module_read_master_readdata -> crypto_module:avm_read_master_readdata
	wire         crypto_module_read_master_waitrequest;                        // mm_interconnect_0:crypto_module_read_master_waitrequest -> crypto_module:avm_read_master_waitrequest
	wire         crypto_module_read_master_read;                               // crypto_module:avm_read_master_read -> mm_interconnect_0:crypto_module_read_master_read
	wire  [31:0] crypto_module_read_master_address;                            // crypto_module:avm_read_master_address -> mm_interconnect_0:crypto_module_read_master_address
	wire         crypto_module_write_master_waitrequest;                       // mm_interconnect_0:crypto_module_write_master_waitrequest -> crypto_module:avm_write_master_waitrequest
	wire  [31:0] crypto_module_write_master_address;                           // crypto_module:avm_write_master_address -> mm_interconnect_0:crypto_module_write_master_address
	wire         crypto_module_write_master_write;                             // crypto_module:avm_write_master_write -> mm_interconnect_0:crypto_module_write_master_write
	wire  [31:0] crypto_module_write_master_writedata;                         // crypto_module:avm_write_master_writedata -> mm_interconnect_0:crypto_module_write_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [19:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;        // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;         // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_crypto_module_csr_readdata;                 // crypto_module:avs_csr_readdata -> mm_interconnect_0:crypto_module_csr_readdata
	wire   [2:0] mm_interconnect_0_crypto_module_csr_address;                  // mm_interconnect_0:crypto_module_csr_address -> crypto_module:avs_csr_address
	wire         mm_interconnect_0_crypto_module_csr_write;                    // mm_interconnect_0:crypto_module_csr_write -> crypto_module:avs_csr_write
	wire  [31:0] mm_interconnect_0_crypto_module_csr_writedata;                // mm_interconnect_0:crypto_module_csr_writedata -> crypto_module:avs_csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_instruction_memory_s1_chipselect;           // mm_interconnect_0:instruction_memory_s1_chipselect -> instruction_memory:chipselect
	wire  [31:0] mm_interconnect_0_instruction_memory_s1_readdata;             // instruction_memory:readdata -> mm_interconnect_0:instruction_memory_s1_readdata
	wire  [15:0] mm_interconnect_0_instruction_memory_s1_address;              // mm_interconnect_0:instruction_memory_s1_address -> instruction_memory:address
	wire   [3:0] mm_interconnect_0_instruction_memory_s1_byteenable;           // mm_interconnect_0:instruction_memory_s1_byteenable -> instruction_memory:byteenable
	wire         mm_interconnect_0_instruction_memory_s1_write;                // mm_interconnect_0:instruction_memory_s1_write -> instruction_memory:write
	wire  [31:0] mm_interconnect_0_instruction_memory_s1_writedata;            // mm_interconnect_0:instruction_memory_s1_writedata -> instruction_memory:writedata
	wire         mm_interconnect_0_instruction_memory_s1_clken;                // mm_interconnect_0:instruction_memory_s1_clken -> instruction_memory:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                      // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                        // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [3:0] mm_interconnect_0_timer_0_s1_address;                         // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                           // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                       // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_stack_heap_s1_chipselect;                   // mm_interconnect_0:stack_heap_s1_chipselect -> stack_heap:chipselect
	wire  [31:0] mm_interconnect_0_stack_heap_s1_readdata;                     // stack_heap:readdata -> mm_interconnect_0:stack_heap_s1_readdata
	wire  [11:0] mm_interconnect_0_stack_heap_s1_address;                      // mm_interconnect_0:stack_heap_s1_address -> stack_heap:address
	wire   [3:0] mm_interconnect_0_stack_heap_s1_byteenable;                   // mm_interconnect_0:stack_heap_s1_byteenable -> stack_heap:byteenable
	wire         mm_interconnect_0_stack_heap_s1_write;                        // mm_interconnect_0:stack_heap_s1_write -> stack_heap:write
	wire  [31:0] mm_interconnect_0_stack_heap_s1_writedata;                    // mm_interconnect_0:stack_heap_s1_writedata -> stack_heap:writedata
	wire         mm_interconnect_0_stack_heap_s1_clken;                        // mm_interconnect_0:stack_heap_s1_clken -> stack_heap:clken
	wire         mm_interconnect_0_incoming_memory_s1_chipselect;              // mm_interconnect_0:incoming_memory_s1_chipselect -> incoming_memory:chipselect
	wire  [31:0] mm_interconnect_0_incoming_memory_s1_readdata;                // incoming_memory:readdata -> mm_interconnect_0:incoming_memory_s1_readdata
	wire  [11:0] mm_interconnect_0_incoming_memory_s1_address;                 // mm_interconnect_0:incoming_memory_s1_address -> incoming_memory:address
	wire   [3:0] mm_interconnect_0_incoming_memory_s1_byteenable;              // mm_interconnect_0:incoming_memory_s1_byteenable -> incoming_memory:byteenable
	wire         mm_interconnect_0_incoming_memory_s1_write;                   // mm_interconnect_0:incoming_memory_s1_write -> incoming_memory:write
	wire  [31:0] mm_interconnect_0_incoming_memory_s1_writedata;               // mm_interconnect_0:incoming_memory_s1_writedata -> incoming_memory:writedata
	wire         mm_interconnect_0_incoming_memory_s1_clken;                   // mm_interconnect_0:incoming_memory_s1_clken -> incoming_memory:clken
	wire         mm_interconnect_0_outgoing_memory_s1_chipselect;              // mm_interconnect_0:outgoing_memory_s1_chipselect -> outgoing_memory:chipselect
	wire  [31:0] mm_interconnect_0_outgoing_memory_s1_readdata;                // outgoing_memory:readdata -> mm_interconnect_0:outgoing_memory_s1_readdata
	wire  [11:0] mm_interconnect_0_outgoing_memory_s1_address;                 // mm_interconnect_0:outgoing_memory_s1_address -> outgoing_memory:address
	wire   [3:0] mm_interconnect_0_outgoing_memory_s1_byteenable;              // mm_interconnect_0:outgoing_memory_s1_byteenable -> outgoing_memory:byteenable
	wire         mm_interconnect_0_outgoing_memory_s1_write;                   // mm_interconnect_0:outgoing_memory_s1_write -> outgoing_memory:write
	wire  [31:0] mm_interconnect_0_outgoing_memory_s1_writedata;               // mm_interconnect_0:outgoing_memory_s1_writedata -> outgoing_memory:writedata
	wire         mm_interconnect_0_outgoing_memory_s1_clken;                   // mm_interconnect_0:outgoing_memory_s1_clken -> outgoing_memory:clken
	wire         mm_interconnect_0_timestamp_timer_s1_chipselect;              // mm_interconnect_0:timestamp_timer_s1_chipselect -> timestamp_timer:chipselect
	wire  [15:0] mm_interconnect_0_timestamp_timer_s1_readdata;                // timestamp_timer:readdata -> mm_interconnect_0:timestamp_timer_s1_readdata
	wire   [3:0] mm_interconnect_0_timestamp_timer_s1_address;                 // mm_interconnect_0:timestamp_timer_s1_address -> timestamp_timer:address
	wire         mm_interconnect_0_timestamp_timer_s1_write;                   // mm_interconnect_0:timestamp_timer_s1_write -> timestamp_timer:write_n
	wire  [15:0] mm_interconnect_0_timestamp_timer_s1_writedata;               // mm_interconnect_0:timestamp_timer_s1_writedata -> timestamp_timer:writedata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // timestamp_timer:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [crypto_module:csi_clock_reset, incoming_memory:reset, instruction_memory:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, outgoing_memory:reset, rst_translator:in_reset, stack_heap:reset, sysid_qsys_0:reset_n, timer_0:reset_n, timestamp_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [incoming_memory:reset_req, instruction_memory:reset_req, nios2_qsys_0:reset_req, outgoing_memory:reset_req, rst_translator:reset_req_in, stack_heap:reset_req]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	ted_crypto crypto_module (
		.csi_clock_clk                (clk_clk),                                       //        clock.clk
		.csi_clock_reset              (rst_controller_reset_out_reset),                //  clock_reset.reset
		.avm_read_master_read         (crypto_module_read_master_read),                //  read_master.read
		.avm_read_master_address      (crypto_module_read_master_address),             //             .address
		.avm_read_master_readdata     (crypto_module_read_master_readdata),            //             .readdata
		.avm_read_master_waitrequest  (crypto_module_read_master_waitrequest),         //             .waitrequest
		.avm_write_master_write       (crypto_module_write_master_write),              // write_master.write
		.avm_write_master_address     (crypto_module_write_master_address),            //             .address
		.avm_write_master_writedata   (crypto_module_write_master_writedata),          //             .writedata
		.avm_write_master_waitrequest (crypto_module_write_master_waitrequest),        //             .waitrequest
		.avs_csr_address              (mm_interconnect_0_crypto_module_csr_address),   //          csr.address
		.avs_csr_readdata             (mm_interconnect_0_crypto_module_csr_readdata),  //             .readdata
		.avs_csr_write                (mm_interconnect_0_crypto_module_csr_write),     //             .write
		.avs_csr_writedata            (mm_interconnect_0_crypto_module_csr_writedata)  //             .writedata
	);

	crypto_test_incoming_memory incoming_memory (
		.clk        (clk_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_incoming_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_incoming_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_incoming_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_incoming_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_incoming_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_incoming_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_incoming_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)               //       .reset_req
	);

	crypto_test_instruction_memory instruction_memory (
		.clk        (clk_clk),                                            //   clk1.clk
		.address    (mm_interconnect_0_instruction_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_instruction_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_instruction_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_instruction_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_instruction_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_instruction_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_instruction_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                     // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                  //       .reset_req
	);

	crypto_test_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	crypto_test_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	crypto_test_outgoing_memory outgoing_memory (
		.clk        (clk_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_outgoing_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_outgoing_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_outgoing_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_outgoing_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_outgoing_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_outgoing_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_outgoing_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)               //       .reset_req
	);

	crypto_test_stack_heap stack_heap (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_stack_heap_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_stack_heap_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_stack_heap_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_stack_heap_s1_write),      //       .write
		.readdata   (mm_interconnect_0_stack_heap_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_stack_heap_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_stack_heap_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	crypto_test_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	crypto_test_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	crypto_test_timestamp_timer timestamp_timer (
		.clk        (clk_clk),                                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 // reset.reset_n
		.address    (mm_interconnect_0_timestamp_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timestamp_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timestamp_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timestamp_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timestamp_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                         //   irq.irq
	);

	crypto_test_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                      (clk_clk),                                                      //                                    clk_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.crypto_module_read_master_address                (crypto_module_read_master_address),                            //                  crypto_module_read_master.address
		.crypto_module_read_master_waitrequest            (crypto_module_read_master_waitrequest),                        //                                           .waitrequest
		.crypto_module_read_master_read                   (crypto_module_read_master_read),                               //                                           .read
		.crypto_module_read_master_readdata               (crypto_module_read_master_readdata),                           //                                           .readdata
		.crypto_module_write_master_address               (crypto_module_write_master_address),                           //                 crypto_module_write_master.address
		.crypto_module_write_master_waitrequest           (crypto_module_write_master_waitrequest),                       //                                           .waitrequest
		.crypto_module_write_master_write                 (crypto_module_write_master_write),                             //                                           .write
		.crypto_module_write_master_writedata             (crypto_module_write_master_writedata),                         //                                           .writedata
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.crypto_module_csr_address                        (mm_interconnect_0_crypto_module_csr_address),                  //                          crypto_module_csr.address
		.crypto_module_csr_write                          (mm_interconnect_0_crypto_module_csr_write),                    //                                           .write
		.crypto_module_csr_readdata                       (mm_interconnect_0_crypto_module_csr_readdata),                 //                                           .readdata
		.crypto_module_csr_writedata                      (mm_interconnect_0_crypto_module_csr_writedata),                //                                           .writedata
		.incoming_memory_s1_address                       (mm_interconnect_0_incoming_memory_s1_address),                 //                         incoming_memory_s1.address
		.incoming_memory_s1_write                         (mm_interconnect_0_incoming_memory_s1_write),                   //                                           .write
		.incoming_memory_s1_readdata                      (mm_interconnect_0_incoming_memory_s1_readdata),                //                                           .readdata
		.incoming_memory_s1_writedata                     (mm_interconnect_0_incoming_memory_s1_writedata),               //                                           .writedata
		.incoming_memory_s1_byteenable                    (mm_interconnect_0_incoming_memory_s1_byteenable),              //                                           .byteenable
		.incoming_memory_s1_chipselect                    (mm_interconnect_0_incoming_memory_s1_chipselect),              //                                           .chipselect
		.incoming_memory_s1_clken                         (mm_interconnect_0_incoming_memory_s1_clken),                   //                                           .clken
		.instruction_memory_s1_address                    (mm_interconnect_0_instruction_memory_s1_address),              //                      instruction_memory_s1.address
		.instruction_memory_s1_write                      (mm_interconnect_0_instruction_memory_s1_write),                //                                           .write
		.instruction_memory_s1_readdata                   (mm_interconnect_0_instruction_memory_s1_readdata),             //                                           .readdata
		.instruction_memory_s1_writedata                  (mm_interconnect_0_instruction_memory_s1_writedata),            //                                           .writedata
		.instruction_memory_s1_byteenable                 (mm_interconnect_0_instruction_memory_s1_byteenable),           //                                           .byteenable
		.instruction_memory_s1_chipselect                 (mm_interconnect_0_instruction_memory_s1_chipselect),           //                                           .chipselect
		.instruction_memory_s1_clken                      (mm_interconnect_0_instruction_memory_s1_clken),                //                                           .clken
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.outgoing_memory_s1_address                       (mm_interconnect_0_outgoing_memory_s1_address),                 //                         outgoing_memory_s1.address
		.outgoing_memory_s1_write                         (mm_interconnect_0_outgoing_memory_s1_write),                   //                                           .write
		.outgoing_memory_s1_readdata                      (mm_interconnect_0_outgoing_memory_s1_readdata),                //                                           .readdata
		.outgoing_memory_s1_writedata                     (mm_interconnect_0_outgoing_memory_s1_writedata),               //                                           .writedata
		.outgoing_memory_s1_byteenable                    (mm_interconnect_0_outgoing_memory_s1_byteenable),              //                                           .byteenable
		.outgoing_memory_s1_chipselect                    (mm_interconnect_0_outgoing_memory_s1_chipselect),              //                                           .chipselect
		.outgoing_memory_s1_clken                         (mm_interconnect_0_outgoing_memory_s1_clken),                   //                                           .clken
		.stack_heap_s1_address                            (mm_interconnect_0_stack_heap_s1_address),                      //                              stack_heap_s1.address
		.stack_heap_s1_write                              (mm_interconnect_0_stack_heap_s1_write),                        //                                           .write
		.stack_heap_s1_readdata                           (mm_interconnect_0_stack_heap_s1_readdata),                     //                                           .readdata
		.stack_heap_s1_writedata                          (mm_interconnect_0_stack_heap_s1_writedata),                    //                                           .writedata
		.stack_heap_s1_byteenable                         (mm_interconnect_0_stack_heap_s1_byteenable),                   //                                           .byteenable
		.stack_heap_s1_chipselect                         (mm_interconnect_0_stack_heap_s1_chipselect),                   //                                           .chipselect
		.stack_heap_s1_clken                              (mm_interconnect_0_stack_heap_s1_clken),                        //                                           .clken
		.sysid_qsys_0_control_slave_address               (mm_interconnect_0_sysid_qsys_0_control_slave_address),         //                 sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata              (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),        //                                           .readdata
		.timer_0_s1_address                               (mm_interconnect_0_timer_0_s1_address),                         //                                 timer_0_s1.address
		.timer_0_s1_write                                 (mm_interconnect_0_timer_0_s1_write),                           //                                           .write
		.timer_0_s1_readdata                              (mm_interconnect_0_timer_0_s1_readdata),                        //                                           .readdata
		.timer_0_s1_writedata                             (mm_interconnect_0_timer_0_s1_writedata),                       //                                           .writedata
		.timer_0_s1_chipselect                            (mm_interconnect_0_timer_0_s1_chipselect),                      //                                           .chipselect
		.timestamp_timer_s1_address                       (mm_interconnect_0_timestamp_timer_s1_address),                 //                         timestamp_timer_s1.address
		.timestamp_timer_s1_write                         (mm_interconnect_0_timestamp_timer_s1_write),                   //                                           .write
		.timestamp_timer_s1_readdata                      (mm_interconnect_0_timestamp_timer_s1_readdata),                //                                           .readdata
		.timestamp_timer_s1_writedata                     (mm_interconnect_0_timestamp_timer_s1_writedata),               //                                           .writedata
		.timestamp_timer_s1_chipselect                    (mm_interconnect_0_timestamp_timer_s1_chipselect)               //                                           .chipselect
	);

	crypto_test_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
