// (C) 2001-2015 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
H6QpZOH4BZoNzN0TUlNkDK1rHlFyQWV4lPu9JD987PgVHNYO4nO3R9wRsXIxXkqljOV6Zh2pDKdc
FtzAEgGbta6P9HIDq83gFwj+tRHh7HT362bQ0bhodsJiAUxC0/BT43WcHZPo0tUsA+V2RNij6JjS
bzk8tQgsdaqx0w3t0SZW3L7MWxy00QRghScb9WP14ajjGZWr6BNOqsYRSNlaFGY5El6W9KkKnvWP
v+DQXMSV2SyZ+pjPKuL+j9lXFQmk7jD2wlQDMBsbCQmcNexrFzdO80G/mDDY2Ce2Uh+JzW9ijZ0y
Q+jtwxXA+UCYH1tPHp3hYIoK0BLV9eSDlVj3pw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
uqFo4QPAqfimJbWwNsEhCb6Di/ZABydrfOIPFcqxs5Fuaih1TdttabgvKqrxy90kNYCqwAnqfU8c
PgmeQ+vw+MbQR3NRj8Kwd1bYUVKbhNcKw7Xc65I9XaQXpyazTxjJ0o7dtCq+fLEJ6CcmtMOwk+S+
b8CH//Kni388yHla45sjPownsbRYk+QAz/2WdWbV3gxMaqftjjdOHJSAE9X8Y2AYi0ehsCXZjIUl
2rB/ilUb7QGjGkqi59sU5p2w9rRDwDMSk7tdrUfdgrH3R+K3KayOXPdRElQj/am41x3Wjr56iqIG
rwRRFQk2/jifV4X4ciGBYfZZuLWjdo/Y266t1WE7AvBRPn/kpoWi63usD64H6Dm5stYhXj0AwzkV
xSUA0Wy0hJpK6//WUn7kA166XMvg4yLrYBmmTCUWA0H8GD9uyYtu3gBOuYie8ZUYHp/4fMXjP2Fq
rksbPcOZlUQlNqXaGlO9qfZ+IbLOLqtc5hiWGWHF6lohj3Nlb4ahMH6YXyR0AT3oGX+DwPJwc7Ek
rR70tIekV91r4eMkhx7iTVZsxyEJqGBIplaiul3PMvFzPeH09N1S4Cu6ZyAbNa9nDht+bJyaY0NB
52bn+7BTkMBov0HT4lLSTvQz1Im3px4M2pm8LwaawIAXboyfCX12OPMvRqXd7Nf2s2dZ8sA6xcne
pmQR2/zfbaOSN/Xe/PLHo3nOivbOjsIlHVNZHOE7efAuEaFL+UhcHCRpUEz8B+6qp+M8ecHHsfco
0+DJVutdLGOs6cH9nAKNkPsfIbGYO/Y0Rpf+Bpj2tVNjB7XlupyyzSsxXuTO8arBIt1KZIPwdUa2
pTZSY9BEQ45L8Aii4bOZ+hhJ02CtTbAQroCoRpnw5hI/sOipYNNDTli4njuj67pSM5h1wubp2Qr4
k+2E1YQUhDAm51DF6hhAo4G+Fwkoc7u44yarKgzhYfDjWUHP+kfwpL2rLEJB+Or+DZ5o8RcNWMZg
3Q0Y/LyP4/eFWBxwFnSm99GfTMBaaJYR90G/sYmGssdOHV0zUKclj3mruBhVbiYvaR5YO1UQbTBt
yrMRQp0q/Kjs8HBTXvwjnCET6dfqLiWvkobrYCBuUW2fpTl1IZNkRp1Aq9W/RXYXzOO/cg6M94k1
3ISiPH2F0nwGYXfBNVxoREA14O5bv8UQloWYS8cLmdrkgMI2LDf0YVrVYkhKB06j/ddfqk4PTPDG
XJCQszRiu6MQ41eqPoG4/wonzPPfb2ly6ZpyMEUF8Oq0KZ3Ow6OlpXcwKzCiGU3h2gD9wxzCxD9Z
UM9+S4kW9hwKXTcoDCghBUgtwLFlTkSvma+/57/K7yDJpT7dPGtyepcI0i+pW1+8UmuIXLxsAGK4
HGY6Cdx2Nnue9z+2Q0VLrC6250u+HZn2r6goSSiyA0JWjbV4J+Vjnpb4suXKD/0P58Y45UB+lArc
zr1V72cmKZ9z1lqvDM36nE1zVmYEI811a5tnEHWht/0xJnIoCoixRANBjTW6m+8NBi6r+aCoeM/4
R0I1cN+ktqnnEWXj27O7USjdM82aEsuWfrgTeri1XdSzcSD/gXPFz9tCEAjbi/F1HuMrgb4joN6M
rAU4PvS4+afxsxo/C3aMkmgk8vf5BwsEdWtip64RAarDDSiUyhlJs8uf/JlY6zjbc3AMPj2nVxQ7
p8uFMyeP8ksdb/kkYOf99VfXC8aLRlhXL64eN12Xb/0XOK6yyW9rH/EIU7/GgusexugchOudaAGl
H55YdCiximsJ5KF5r9Bxjt2z7Zx2sRJA0yltMJnc6CzlJBWfvB0DsZnKb4rpZGujg+x3DJ7rg06V
0UUeB2U8PMMu2IcYBbRfF16tgQI2uRmt1yZHq25ZZE1yJieIwoNqNRoQUoJJ0aDnhFjQjB7+5xP/
uFj7SXKCDPLtJgzwBPjbRuMuyYkhQH6T98zt7jnl7PSTlpUoJlGbJW2JqtSQC7RY3eG8z8gmD5J3
oueIFkchbvIiSamgwx8xGvhPrHcTUAptt+d49EqnoId7bNJCw8Hutl4EvFnDvVj4lMafrh+r39yS
coCFRHctB9DCYZqYilz0F3XnfOyQ6cINM2BVLxbsFnE0w2YJdqKVt3RSGE6u8HrlkAL5OsyZuQa5
cUoxIW5GJJEnEn8d8k8b3/GjLRu8XmTyDBOISVIxehUpDF4BzphzJcDideBGI5imlGespyqRvoPY
rU2Br2IiB5HForKMYtWqvj1cqkGzTZfEsseo0bFkqaTYBqFPV1AC7PcY2sUNPPkL0j2muWMj29wb
qRhD6uN8Lba/R7GJkicIPFuqfcK71841cwCgYsoKImFF6+Y8nJTVvF7rAKKjky792btr0OFJ/cTz
dRKr6zbDDOzoxD95+P76fGfbF0y5UgAuKkfFLGvUtyL9uKzkILyGq9gktjRkGVR9ErlxGh4gNnXR
WENqw3M++hWZojX01kNxG2xGMFgVej47tAAwNasz5NyqC/oYHU/Zzspe+s/gCzdupF+PjpI0gPKj
tZcL6bpzFdyrxjRjffL8WYr6dpepbKxFOgTx18yyt/lrZBKUXn5ybF46XiWqnBd75f6nV6Wreoao
9masF1gUvxGPyFQW6Ruu3zLBHmZ17sGUM6Bzj9kCHdI7DLygkq8TpSr0jvliLTJsKidNSbG9rqSb
4Cbbnxsbsvmcs9Lsd25bYfav8SYR5LOYIJQ/GvHjGHTE2fs61eLp9axWQVDBPqHsXFSR7UmKAfgr
hf0nynw9WGZXfkJLYTq+L8laiZxENIcNWhRogv3vyD0RSD18lj4+Atub8h5/wfE8Sj0wNYyY13Mv
AXhXHjvN1iY6w30fqd4MLaH+liT4Qqvu7dOPtRoQzJIKEQp+uTOZPlES4vUhYWJO9PQpBBIuYSfK
49CspdJgz/L4SUAaEuMZOmiaZx08nXhyOzmFq0SG+vLuK5/RcM+KCs4SjvktlnU2SsRwA6xcjo98
JxIyjsJkKRTULjwNMv5QQMPyWcQpkOETdSbDQw1mW8OFGB27SZqyXra5mUxzot7WoLFxdKvj/8Z0
k5PScUO2+0GJe7Cp0uPMGGpQbaFt2MBHFQClOP8Gsjkr9coq8QS9mWK5GxoqPPtj8UNg6O9J7UyF
tfgtySe4K2yxyW0M4GcJ5RNECMOQfDwX552vnCo8xTMGi/eJgGHtyHc1ZaGWrMsYXTjcuzKJa3Dr
DNTb0O7F9IOucgsnNuEqrMxYDEZDtuWFfoellwd0cSXXhJmaaVLB+iVk+c/X1pJqku93RDIesMyE
8GukCe3dTan2p+kylQNf0AxYOIjr3A5/3TfiAzVLP3dg1cY4EoFrg7/iZpkU2j1EGx1K2iOrrxo/
PHVLogQ/fQ2BL4Ix1ei9+7s7K8drY3V+DFwoayUgwuhzJIOzKmzH61wcaRVp6NK7f2wkU7PMlEAO
19OS6/JNnQNqRSO3wtNOOF5BMmQNA5JZiWRioKvZ+PMFJ/MoOOwHyMI2fW7Y3Tj5stYE2QMzu3b0
eoHUkSwy81mccvH/HmL9w9lBiykG6I639z/NJRY7+LLzcNvRsQvIV06YoR0Mqk5NjZQn531/FF9Q
NDH/jZ0y2iUjRB9Ori6yKrRpvRctujjjqtMdcrO7iH3GPxd1QLTJkyES6pEeQx8FsvYnVfVuvX51
WqktrqfU4xnhr8LfEEq8DrypzR/s75ZDHjsPHi8StkhljIKa/Gf0UR7c7dy979SxSBJHQ77G8l+k
JAcAVxtX0OocotWpwTXUmeXhTkQ039IDeacOXl7ooPfCS8IGGjGXSo5i+VfpU7eJ00YOTPt31fwu
HXGoz6G+nWoPzHBqqZNqwZlEVm6+FGAIiHevxJVQwYD7+M69776ZgQ9+OQnGddJpXlriqyaDlNTu
wJzrB/AIpaF/viF4uQog0pGdTTo8eDehga1W5GGWwZCyldHs5ys4Ib8v5DBtvSGkkhpaXwlS752d
tizEjZqRAIpcrJ84sOiZmPd5cPQjIyczA2egiGBD0/bSeEymCys5A+eD3haAVAdDwqqMW5Uyrhrs
B05/hENyD8rr2A0FwjmWt2zLCMfvfB60x5kGHXfERBSP19GlRBplC757N4Vv6NS1IqrwpFNl21Ld
w1SlQ5NJTkWxZYLhe4lkT5Kekb1VKxGWFEA7yiYDC92oAoAs9P1+4wPYfdrCk/CEIySMfxYBQy5x
7ZghckHBsFepAp7pC1+r+j0crNEBkHgM5hvp3DEmJZqXuD4mDE0FAwy9Ju1fhyGGixk2cJ2ql3lt
6psULb6KRv4ECuSo/V/QFRFKFP6fZbe3O881KcB4DWAsN4xGkI/tHAGfhCDUjaUr5fgyAYZxuewV
HrZO49JwqOPEweoOF9lEQTpE29qU0AmgxiPE0k3eKHMjRyandogs+gSGETlNqsxX5SrfEN8J1yd8
YfFnaEJpWE0+osATeULNVqkI0OHe1mV+QttQLofRoAy6v/zlUUHgjo5efqgwphvmz9Jnc4yGzHpH
s0RF2SIckVap9wq7PRwNqJbblk+mwHVKb3ZMCWV2uYIi7uMcecOtv+ziQxbvXDXuM3sGRkV+mv4y
WzUoyZdBxVfQv5okOqDdLB7yxZ6In7Rd0Ygje39dgX42gu8lG7UZuOf/SWXZlbWLXHd3Gwmvh6mg
n52VnVmug9MQPdD+/lRSI/I4lPaXzstF+g0jMu7SVRoLg7BM/iku+qp7GIH4Fx/keMqydiNyHmlS
KoBvOsVAgx/W547VcwfyZfd1I3jDziqk4AjEHqSxEUDTTj0NZL6SqK9Y6nuoiX5OLAzciVEw/CH9
HSGSlB16v8CkG7FlsI6aMGvIoiZE+w0OPQu4v30EBgacWFE99QtW4BFyW0BuDe0qXW3rz5CIFHxd
cUnBPrbF7uLsuWR3kVzzzhewroTXS/SWm6iZ7SSAv+PfTxL2l1mWm+e+XADCUIg0al+/G+zktmJi
Nr7NbdS3rCOS+qIV2Afai6Fs37Jp49mJszfB6evpMKFKmSnv4I5ZvI0j+6Qfph/jxquu4543AfpX
BiiJasWYUpZkl7ZvBDtcMvSH4ULhiHaJfL3k3cg+LgD9RWi9oT2ykujs1CylMUIWrrHWtkcnsy4i
JJsqd5ym0yegh2now0DpzmOVj6TrmlrbQpzlO0Qx5NOC86WvrYygEpyAMUPK0WTDlkDTWbCkUXN0
5RLnbqEKex8mWLPq485hfmtd6PPfuj5/f4cvJAu/RgrvJAwh1q48HZRgrTQmWkPFooEHieuKllXk
U0Pb2VaN3LQzMNdTMh8t0LzLbu/s4YQb+FcBvvPYwxUcchDNTPbKWLcXeuFqnmN8ttxSZAimJVQY
T5M3N+x1LD6V9MzkxCANf3yBeE+acVNAbqWoMEX2phEaytI93Mgq1lSZTBKhr3j5RWwEMIXis6eE
cRQXASCOE64WODkcmOXCxE76g0o0PomWmN7jsYLHGgU9rBLKJxYS9l4KykiAlGJjwTwOkt2vE+gk
OgL2Yfj0UzJEGwkEHSlQRPUqSeF8QW2ZFc68iOKvnDTKf+7Yr0+kjYul7FBQxR5MDGQQNJ2xtn5A
Dfjq4Y5aHaiWpvnkD0If3j0FrTPBMrvlaUoMATH6n4+5UNq8qOjfxj+JEcdXr9BEnLSl2aYJDOx/
i7OPVzZZZHiXP4gFsEEsK1DcCs558dSsJuzi9h8chyXF+pQ5o6IGOAj2r92ElQSz3y2Ee2Xt8S9J
WdcDHGTJldr7IyaWeLNnhvOwQXuQka6J8BtTpVKfyURLQv3khlDJV1o13o7OlplGvscMnUfxk3LW
Ogxu9TV8J1KkwPtn9Os02P8/TiNa6IHl9VQ48I6LTN2PTAh8M5DXPB91GmEX/QM0m8yyI/l7v1aB
2fcEJD1lkiyDCj4n8NslP2aURoDM9smXpAVD/I/S0AW85ZXCMByr8KKE4bxO1nSxA/UYgbgXcQK0
Xi7P9ddUIUESwSshgCtVqMrePLTQcgJj6nCdax/gXIe0wQcr3odZ7b89LlBi/O4pkR7cLG58yWaB
SukTMn0zGqx2jO4Jyp3PskZQLAvy7P++h3CmbEbqteaJldO5Kg76qg6W1I1kqRdlFv4SUGb1APK9
cmKThEyqnsGxSKSdLkT/1tFiJaBYfZxJlGzhEKwY0rFMPC6U1BW2C+CMpVo505er9hBkq5VQ9eWs
nDUVypSAJSwdy3ZNvEvX0LgmPXAYHJrDoaIA4n4Y6JWZ1N/OGP2cjA4QbytiIOB24Fq7+eMfOKyO
maEg5QaBfYwghGWqGORNfJrH3iHStFGFpKJ+cvr/IgMHAIs6CeuNrnSL7uO4ORAY4lVsFSo6WWSG
IMK+CU2cDD+u6Jz4Z1Yif4qrgooo/ZWKjtd6GA+RfHRhWgwhWFLEGePHx+85lRs/c7+FD2TMgdDI
AIJ7IZ9RhFjKAXBUDnQZX2cAmCSfHBUHQqDP0DHYx8RbplB+BkkAujEcpnMzQDqZbJdjgqi1VWc/
SSOVa8Pq0rpJjD8oSwHicJEWuZYKjvnXil7bsI2lzzNZL2kfvFStJTPmtiSC/UU47wTAJlkSZOkQ
UU2xymxAuKIcDyt4ITPDVLnM14wssS0Yx3ivYqxeDxO3Lat15V0k91JW6sCV4xHD+1TLWJlZca8P
U09XCvgSe++b7e7iSqqpEiQjEDiheDYBuLi6nUI3iVuuQIzUgW4bSW5J6YH6HCo4UYJ9GXKlooU+
LN3LR6lSb+Ir0Hg7FtXTerwZxG8re8t6p1RjjeYaVYdcEJaDCEzYQhlEOMrFI++IsZr3+LqNTmwG
56ZYzeC+cTIB0fT7UWCKIjnCJDCzSFU+o8JUMr3tzROrUY+Gwtn/vzSB8fcAndweyryM5Nht2FsA
t2uw+JyWBdm8NRVl4NjH8Oyycf4IT1GF/Oi5Tgd5nnipZDOkwNuFFCasA0h77HLOF87eN7s0Bv1w
f/KQAt+nfcE4DGUw1o238dMW8Rmng06wsis9zc3NA26IYs5C9s26fdE60uSGuBbnGJBxNbjRD+p3
dqr/UsUnEzaT01YRM98lagtjoLyH4JPq9/TqNkb8NrmD9j0JpewrkdqDL3hKhIDJIDHFCX2qIg2N
om/Z+5Km9L5ygI6y/kO+YVhOTlfkrB/DE19luPSvVPYRUADt5+nBKVzP0DUNEFLGQiBdlxTV1/w7
o/ZNGhXu2aa4Q3suR+EDQmsnKU+hzNQzwF5ILo7IoCk3xYh3xWVWjTVsnAJBMrraqeOhj9Nu/Aau
aqwz46/jMUdv+n6yAwO/FS4dnAtsgpNRXLpGE3gxhknh0cSkWoggoIb9yCE0y5wMu0kA52RRliJg
4d3Ljp4GvCTlxKX8f83i8xhqoCsqg5QdCtd8GE5mCqWDQOZ9WKklGR5KXHtyoi4zfE4T/cruKVe4
PsHb+a+ATex5l2FH9Z515Z0iH2KHuZmCik/0sRu4xqeAP2yQGeRmMymPAL4KUOILJB9yPRJBtBN7
rwVonPLUVkUPIit936omxN7Hk/CBERWA4ehXVb5Jv2FwYE34kRB8U6u4PEYrO+vbCCw2EKf3Aw0L
fRcOwo+88/BctWOWYCXrJAT8ncQUVCnDmFFmsStI5KMOq0j93DTE66MIJXeDvatVczLaEc2RaSve
/19JoxExWRCpUBfu7Ud9UnlIOxJO84hX81i7bAQumd14Nw5rs3k7IpkCWPrT8suqIScpLGsq1Lrb
AVtuzJ4dguRSTZD+C/hDoR6g39CHCujO0zhV5b6H7lmvWmHGi9KXpQEnfYcJ+p2KXC85QH+P7pe8
qOiV93WbLGpeca8WRbrjOYRo2JUx/VtGqZ9F3M/SXtwqZ94FOoUDZdPFl4DE91/TrDb9aHjX+SO7
UX+/lsqofdmRZ+wl/R9LSjphVSZHG/kqatqcRyW+rw+9Ir7eH4MrXLZ168kk4tp2qqr+lRT+hxyT
V8Xbf7VI5e2HCgAoYdmSENdtlQpeJhSvHBUUMDhX4lQmbYnxuI3d/QgQ0T0eiCCjdtEyOIbeSczc
Nk012LH/jjLi2nQxx+xjVRY/dFuUhpMjWP+lLz6fach1IttmbRBUWf5Gl3fckyYI5JkAK5JYBZHY
ltQlfwoR+cR8t/DzBuxsnCg8YTcpFLVbTfGs9427gz98kjS8vTylYPe/BuWuv0tItw5E+1qQ3ZDj
W76lm5Ew0RfudNW0NkmqArwKZHvYPSms0hWXrW6vwJKe6LRF1fBJ/3KsqI/F7elevDj/rmKa4xuw
jkvfnXrEYG+sHePfZ24O1682pc2LdQNAUxNZcGH7No64hP+6JQ9WJB7GjlBGc2OLeNY1ateZF/ej
U7QUEDiGrCe+cqo/57pMH9o+wuoKNXWY5KlkJmXYQhwCVH+zRU/g3XgU/uOlm3mlWPJ1SiltykGK
dhVhvRWLe5DPz2vNA1IX2RyJMf7Po1H8/OuVU8GE7WOTbZ96VwkBx9NdGtuUVzpaqv2jPAl89JYS
oTVkKBQTmMtNjCHepXr0ywflUveTtvkdqY5N02Ey92NuaSK211nyGCqFVw273OLkdyC6sn4VDyo8
Hs5q/UaxFS9jGEOP0tZPJk3CU4exQTkQZJ3AJxC5iHWXkX/5qWzZopx5hYpSpGY62hA4kbCyfrKE
T3yilxZvAbC+Oew8sa8DJsw+IePnig+Z08gXdraZ5jbSrYWU0udqiH+uouVMrF/5FnoRzeKwfT3m
wvaB7CzVkwautLNp18O049o6UnD0x7vUdsr1HeegO3mocwPOcPrKNBD42F4nhF032iHzrgOx2XBU
wBobrNWwxg3kMDSx7PO5Xxk2Dv33j0QzJJ++v3UqAU2BsVtwr1Qk0+JP4ajk36cF0uapB8H/Gi+Q
ML/Qyrnt9BjR1hYePsBemMJPC2JdGvXnfWTJxFczNWn5rra0cqPY6IOY72oQfakaWT1RmOBn0+2B
O8kZG3JBRLLkkOD/63FEl7Kwli9bUMTlYd9VjFWH5nCUIKeYiSIlM6kLIMkpWpSiGJHjJbEqO5QS
/TTMN6jDCMHIcOdOIc5gYQQlKYWJrI8He6OMCHxI7PwOOSOR9EdYSWwU3z6O0HhtfmiXc0cr7VK8
Q1XAhyJBo9lm4Ey2jd7aROGCPgHtiu1xnNPpyzYulD9MjHrEeb+Hw2U2cMqsykPkATnIa0ur3PbQ
fHr2i3GjPXt8F24tj1qe9ltxHqQ4GU9frnChKaGZNi3FGhsfS0rsmgg63QCyn2Wo9GhzlXY8f7Va
BYRBSozbVMyqJQsMB4Xy1NzDlX/Fjhxc3cpTpC7x8h8LM5EH/Q8/bpaUpkCwwWAsSU+PN9sU7h5g
1IttS1MMXBy5c0zkH7Spkkf9pSZdRK9HAzcrwFv2MrBIkvcEqNpI7lJo1xYycMnZqKy+dy4VZUpY
O8RKzjyNbnv9iDvjwBzYZZWwzxTNJu8p8wy9jAdD8E9aO4EyctRL0eZ++3wIS6aFZfagbOE2uL8h
xcWYLyp97s56FQAiohagVNFUhTFMCDk7n6wXiz6NySP3+ehiPKgyablSdaI+Qg9d3PrzA2AdcRQC
WWwEheeTQ0K+zwr9xPD71RVrwP2RGw2w1lQqUit/luKkx6+2RLyIQp8Arl0/9+s0EfO8qqLNwt0O
pWpt2wob6APhvEuKIalDcJJlgipu24KAfqHv0h9jkEtWNED5zGeEe6Kkhd/6ygfNNEaSra9UkDj3
O5mOcg3bk2wYpu+sBQSjLvY7QhYwZ0+sqAtgiA/exWm9YiXwTVqWoAmqOV+THiiaEs1ipfpOAEmP
maKMPzokNv6k8R9ZJPNM8W0QNcwYPvk9eS5J/joKhSXSUHixj6IosdzFv6V4hbE+faIkCHH9+2Q6
Q+4hEm2J6GoAHf2aWQVHAM6G1S0vc/VUncwhoj2tjU1CVjG/B+IjnzC5+i8SPyCtfROIT/e69SXi
MzObad04TRr3L1Buzc+vU3UBda5yPvWvYg5KgqaxyV+spBLfVxWwGNZl54mOBbAuW3g4x1ArOQO8
96e9PlcIbve0EXv/QwQiM+UvMZ82W8QCfScvNInLMuuExIUOgweQ+DzV88+lJXMHhblA9oK3iNSG
HueZPb/ZlbbHuOnjzDodqVEulG2KpK5VljERX/18qGCobPkYxKjxwkpVXtX5kK/EBnvZKYd8vW43
uEyJzeIh5JKw/hSKNV59o/ag1ASH8f3/jpGbg1jZZPjZyIRcdWLKtGaSFIuSY2YZvMcIm8ivhY7D
EZGm3TEEibGgO/F/bb7iEJAFJf6ArME2erIZK21RHh3LXlu/NN/LINGkjPCuP6+7K5WufZpqkQCf
n+ihuHj/30pcHnrTEjxQw2LWtIT3AB1rN8r8WmpTN7Y+tdQc+zNXr97OKsXid9yOBnHH3Il405lY
jE2o4swaEmqPfWIR8VjMzJM9Jq+iALok26Y/FfFwOvd1DXnZKwbWd8m53qEzBX6FnPWNRrtP6nFh
l8yy6w+L50PGhq5mXvT+ePpApZaKyEc6vs1wdT0Ay0aNBUywxRH3CRfaKGUbT8QKUXIvPsHNjQf8
Arr1pTrJXRpAJ6O7hlnm5wnX8mUOzRuN/OafMJ9QPa2k+UbJXCFNGnC0dOU2HZTVOSSmUAATS7+0
UkgJWdfySaJtiwLZhBED8f+6WhwiOBFZa22pP8lxFe06I+q1x3w/OVzYytZ9k11hrPvt5nDsonJA
xCdLrLhyrFz379VB4c7KJ6t3u9N1roIAtd596yEbaZG+Oso1kNmmv3yWXJatIUk0dqYRBGsc6zly
RNvpmavA393KvAe0dWdkqDBMyYtM39PWXwHkuAnq45+gp+5DFHEueJVcU/Ta+rpqbru3o5R7NOrC
xAzWuq9EwqkMrWIhzIRKkygttwp06RFWa2grwea6Jvh5YnAgXfKWijAGSKdblYD+IOTmzK5J4kfN
FfgWvZpQj/X9WtBAR5F6raGDrfgqz8t6ageJsi4tzhZiTah2fsH169Q5BxKnrQy768WF1ztlwzEw
HSxx6AJpn/Fvr334U+bghtsBJjBLj1gsCnkNX62Ju9FNDCPZV+ZTuaz9XIfgzjIEqUJxBfTQzMDK
2PZATQYO7R6+DRTa1NaHJna7bgLcOkhHqATqQkxK1MkKX6IbxpVJUw0R7XdUlWuWk0LmFEHfSyiY
SedJKPAZU1CPRx9Qv0lhnTbZaS1yYM3SZmt2+07eMdkT/xGZ2nF9ylVAh8fxq54chEHQG7nazBgv
NT4170NY/iiThkfMPySXl+6zDJGFcwOJA3n0lC4FZHBlSIARRo6Pjr8WoUkB9kvJNo7AoiQ9rpiC
2g4yV6XSMWXHSuIthqIlbgephmxRC1VJtmz8nWsVouWORzi4ixMtO0X3pZenHBB580Ju8Yp/crDy
YQJNmIdb5Mcn4lPw4pvG1bD1MOtGunY0VD1IUiHrumh0MynFJFz9omWv9vz3vrQcvitkGbSVw50N
f7twfr6eAlrgZS50R/ndK3nVgVAXQ0B24qhu2pGGoxJbO2KaROVLc6zxNXnXTFAKIxaeXLXFKQnc
o27Oq5pbLRwUGEL+l3m2XepMFuoKm0MvZioDH2tt6PAt4IFpTkmC4FLIsV2qd3EZgMQUAGAEJZG0
LBKFD0AEMSG6aLPGFT/MrNnrONb3Q8VlxipfqoV1qAa9WU+BjqWVNSBCV1z+qqjTv39i65Ui7NYf
7pFJ7LZqhh+egOlXequXBvzyy4CT34auwA4u/2CtHrMJCsVNKzgeUiUIm+RWAjjlK4P6IWNK9uJn
Mh7nhdhN1E6p+sZIwB3qRQDqdYPfzYiHl11igJbgDGgpTYbNlkI+HOpaLTQfk4Ga6IsnaKAKYnbl
XFp/JB1j9SV5lC7whJXPccB4XNfB5hM0jgJRB0uy/ZR7KNtVmwvXlP/U6uPZmndqt4XEDmHZ0gBj
K32sRcqRSOYzA6bIzTu4aTdeua7IDp8a9KgEKkS+A4H2RueSMHhknmZfCOdq0eyQfUBT6I1w+lif
xmjxIx87fOpUjePm4xq5Kn8XE63vAb2RGbWF4dEHRi+UlIbRNCU0fJDJNJOdxMjl+z6iAsYDkZZC
xXmkvKg3yg2i+L0+oVJNNN+AnF0xPHQk+gCTHTYp4XP88haDRewTXX/ptt8TCP/mpi04HNq0F25n
Lk5PM+BztlhjpN77IquDqEwBtzUumdr54v5JnbWcyYUAHDZRufWfdS1vrz3Y68Nl08IIb/glWBrM
65bHrFbf1hTWKF9mS31hZsK2taiZdKwmlanqqH7HQ6GRmSs+NkBeChVJj5xkG07TrQXFFmvlUSdA
qovYWalgjKCpnSF0pawsalemgaRQA6w/hCvnWzbr1Ainrj63ieRkowgkLiyHxuOguW6tG5RNjvUz
nEMEGCvh6zSDa4gCSP+m/Yeqmmx35w8hzkUI6ZG2CS/gxwaFsRb3L40QMdCIfnnIHv/oPLRKmsdw
XYLykYa6htbKWNzHLz5BmkFfBBtVw0LR9FAQwKRHcZya330GrSfjL56QYtL7z/G2Y3LHP9ovcnZg
/KBlev3VBHh31yXvgrpXIVTEFR0vAH6Q29seLJaHgN943pqd9hAhy3eSXtqM4dP2t7LZYiZB25pb
x06ZZs5sDO+RcVwlcIUmo1LOJQ420SVOrtw1L00i+KcWqGCmKMq6ulCnBxsr5JL2G/q9tTyBFt8a
WbFk+73Df/0SIaLJSvlPS/XR2Ie40J0kXRsNBzvNWc/8JtdAkj6opKdmZbjbLgsyXafJ9i0lam8K
6ReZYxUZhblQAKjsqJtC3JnfTg+GueTjQoM/MpY5vXNAE/SeMRLePhg/uSZYh6Hr3UAJSgEfpjsb
X1IjXCdEfnJbkshp3KgMQbn3ROYqauQDMEck+I3xU5S9wGjk4iB2gw/4IW2USDW1M400xyhHpjXO
zWyEV7t6rcipfiAq8WNeFQIL+vd+o8RoyTdXvn6O1BabqqYiVc2Kq8j9E2/enEFl3QLnN8sHJRgL
4JuSWkq08e+DMk/ghYltWP0BJhl9O+e+gVkpkU0d9X1SJ/TXUnDvBNTTlgNyRofajuXc1sSnC8xV
YOMxwVeELGSBU0LZwf52tQrxkmILblfegZQkjF1piqnfZt60CnWWrpTXRV9XmTm7Zu+ZXgWnrv4W
HqQCnrhd7mlEbFpJELToZkMCtrOxYXCYQaXyBSWaF4nQZsTAqYEaA4kvOxN3LATQ/SkAlo6iww8r
EH9MFEJeYaxWVz6MmW5G0dn06mqQriBFS8GhLkfdNud8p4rNKJeP8FxjKRsc+tUG0tGzvjeDsbAH
MuQUK/2BmzP2/EwVEYBDGzbZAhELQ5u47eYvpxhS6tlD07duT8WP+G2zP71ehCbPgYh/RYCAfO/h
OnWyISdrLaXbfBBuNgnJuogyCQNHP+NiBgkUQ2uFrRW/xVZeyfae9expFmFV4BGCr+xYT1p02Lfv
J2hbet52aoKvoBLmtvMi0SKdGPLJLmu8QEdrLZ5APCseuz2ozoy1i2parPESmCjO4RQtofe+ZbTQ
+5n5Va6/h9AqgVX5gE8jvJYJKHdjxYa6LsN9z2bz1Qnlpi29sqvPg5r+F2/wQoR4MDHK7NtN/U6X
sXq42NnNCXK1Rgikj11Dj+6acXmMxjIpaBHeKqQGjN87NWEJhn2e5D8or++n5TZryewyEJqtpVHo
whPh6kIcqKYP27aUIriSG6cCokice4AFi7n5J6UHo7UNiwgmsfSyUYGmTzcgLwugYBGaGROOwkZa
TZHUc3s5xzGkeYLrP+O/RfXODYp2hruC+G60uU3r5887YNSriYq4lzhb4PwzR4UQmIruUZAPrSAN
MQXd+tlejMfhEAGM93f8kyl7ekiMH2JVnVeNhrk/FXG+IeUMEqX9QNrwcOsZZLLSFpD0ONFu3aHz
jVGNWT8Um7gwJRkJeNy1A4nsUhTAPWDCYykzd/g3yxQjLRcAfWnMpwIqJm7IdPbUl6tG2TuQSvp+
+km5Glhr941oKRiTXXngDYG6UW0ASci/KbDmxfTEpvfkcpp4Gthgi31M6KCs4fW//aIQ745kITf7
CEEFaAthbpaYkvlMLvmUSZeV3gHspHcvfY383jdzKcycvP69qp+C1f/Zg8puSNljtGi3ye4Fg3mI
MTSYlmuEwNuPaklWNhXWqjsIPoOGmt84xAduzybly7wrSrMZB4FOiuBCMvf8f7x8nYiWEE3/jCBe
Rr7UebTaPUsc6B6EzDyMkGqxNaWjbOF3IIC5twP2yKRKJr+Vpan/DI/L+K6CpeRmML3Mc3J1pQri
yVOfPWX3gkVjiww9K5szum0fACcHb3Vo2WBTnWtJeoKxt9EdwUSgYuHRD+G0AAnpLpNkZRXbq4xu
+/Mlz4uTsu9zmL2EzMwgBoU+D3S8y2fcftsAlYIYIah8XLWBLnlgbe/muFsEQ9YN7U4Qpc2tiaFu
sEJfoRu+KEm8ggtj1nd6/mpfG7I6wuGFp1JnEHcdOX6xBg1j64BwlT16m1z8eLVboXA8027GqTi/
3AJfx4Mx+BBJtubMQ52gf/6lnKi7l0gvBcydZFgZ7Af0goytGt3cePWtRNxRDBeZzLQs+0CITR85
lT50nPiPQVpscKORX9aql0WpBdAnT5Pg2721RWh4UfwpoOZavvxK7VgXHPT8Cg+k2G+y0N4joNA7
EiBDZhT4GCLkkSwWaplMmfptique45WH6lDmGdC+hHPIpfF74955yAF36OU5ZrPuAA3JSxtfXKt7
nc9JT8vsKklAPL/8rw89fdgT8dA9XcYh1FhNZnkyvGvdfmg9ndD/+6BPo8aTxsHjhsPKXQrQ53Fa
gnu/tiyk6MtuOkc2csgaP0KmFiZ3HnngEmVKLBD6DCdvius9vSrcIdsz+oZ5EhlJsf4tKMGa6lHd
/2I0tY2xkNqgBYnt/kfCJSmV0ggTiShj1NK9ZRUwYJnWSwRlL53GY6vo86k+DdJ2afMk/iYBAn60
ZOF2/SyeukiLrRREUWa5vX3311B6zUC0/RwNmidRJCWobFBABz/KZNliv4DVL2MBnhMpf+n5NHlz
miR9Fj9Ihh/UpXCeH3zR+f9sv59AXMfUvsMX9gYYlSxFdAO57BIbIbv1GJMskRkhuW5sT08L+Uaj
BnkJTzyBwoeux/dpd47mCsnFh9ZNve+F4ZxezqxjqJ2Jw0Uej77J0PGqLvPQMdV49Ofth+QUXsBO
TrEN27h3bcn+akPtmDRAhzG5xdVUfpNPCTaTiZ37/lNeMuJL/b8tXUSXVu6L9Rl/7CIg3GchKK8z
FZQ9pW7yporkrOFZbv7PcPjLcWDGlPwEZRVw1x8I5vcqmHN85cR8TPiHbpi/USBcRCVbJcstT+Y5
w8zYz8w5DHBy8qyUd/C6z/eJCMqbnIiac9YJy2UQHykt/dmRtaLnX6IQQyUSPxB7S1oef6PBdmWU
1G3s/dvppMYNONbHRdd9dgzed+hgLBOIEMeiBZ/qNanUjhrx1PbVvhZHUxp+r+55q3amActXtdmt
ItdakmMbW9gGcw8z5cNqISmTVTpCbaxyTclspDtzFnYSwLTYSjLdYFfE+c/qWjkfaDwfKc/UVh8Q
XRAuI7yzvvgAPmaSVbLOm43B7nhvdUP+yXWjlwv17SRl7wnitEPoA8kT2yv2Ey2SIHmSU2m1ZzS7
7+fo72dXX1g8ksIQoETEV0WBEtxN9gB1Shc9QB3jpObx8z9middkNdUVNUxoHQ4sKZtbzWPi/sXm
94FkQ9VnLrVbqnUL1+1mHgImHj97AB9WcEghrZJzh4scLllbCnjOA/Qs4lLSfXVpWKJGZRNrALfY
fBodHgL9oOBYfRlDdZbPG4Gcs1uyaNhLEZeYbqOUjd+qKuXudhUg6uG1zKNZYNRCTwTuyuiU+iiF
HUz7Opn6VQN4YoEDk8yoi9p+DjziYGfUMPoXnp6AFqnKaNTBHOSg/UlvSpQoZdQuvhYb5bPqy3Pt
wL73fpfjZ3rg7p06NYq3qjPosaz8mvOzMPzggKtcKsULnN+6+rbJMho5lnKUEdVR1kTd+WRFV1Ql
heXfevw+xb/Xg4V76xfbXuzabYpNGAcXVpIOAs2f/EP47t27Kd5etQEa4bj7vbN7lHodpjn1u8Fo
fTwQvZSZwNb8o+VR6RK03NPiTMvhe1KZZ+faGLPEn+xtcMb6SZYmzRyxWLmDy6cwoM70T+du9ZUn
+8FPrcEXlo5l6lNXLX4AU3l2XDL0vket3C/WfT7Sw08vfeUokka1QrFERuwZxYQCYiuQT2RsjDma
Fom2wRZPZfWQ65yL57kuvALEkbzueRZExb+D0xcbUIL97iQZssTXn0Elp6+mKY6ASHBNc5v8UoPK
CqQhPHl7DXgwt0m+Xf+3L0SALBf4SV1KufIE818DGy3LLuK7hmmLNWz2IAhPstRD+lhSEn7EseLq
xwlc0Fj+2AxGKswbCV0/ordgZ01cQt151y9JdjNesdqr1G4yWGfs+Fv3tQtH0VJYmHbn3w2Vxz/A
PtxPmX8G0SxwD0KBymEr4boYrv0RMTrMbqWagdihBMRcsNJIXZLJqppjZdWGW0DstM3Uc3LbYjMb
ZpXdKmGm0I9WwI3UzX1GJuBjlpyXeLI4WkC1r9Th9qRpVHtUpZlTSHYwhCNKgeTgZBoOUmJByxHO
YX9B9PiLZyIwCx9icndP6Ad0m9b+tClVVxkL7776/2DRrvh719Omsd0sDWN3odDrJ+cSxok41W5d
cdpKNxXtjc8o9d38QdKysTynqaaZ26wR+IYfAPQTGigt84VBEr6lV7iRm3OySyPlYxM8af55LfOa
B8eWu4/Rv5rPsmtz3UVGl6uC/snvIBqhJXpvX5n1E+8stnyd8YL9icEX/i/YWRJI5SC0lUSSTX+s
/JMl0OH3iNzvZ5k4d30ZGs2mR/cLTdsPWTSX/PBg7lkqzo5FHIls/p/2GWVnwrz5vCsm0EqmNd4n
PPJFZlRSL3d6zNWARHOcyq9LpxBAgcqZfuUAS6XHNJwAUvIjcZkm9iM5B+u1HITdTr2whRtEmky9
BeXq4zYlg32ufBQJSve0iistYhph3OdRPmPjj7T9x7VzQIcvZ1TkE7yavJclpkicGZjbOuNpLf5B
gKSLqv8INuDJYFTZKt9xrgLpG7fiXC320Zc9v1u8nCK6PVUX0xd+aR9V3OathCJeA90EAf80pzFI
LFeCbGNsmDXZ+qKsfPDATzDVBjhIBxJ1DnsQOxzpIGZqGakHROSl+V8NHTpqUdfs7nU9PkzfdR33
C87i9MNwy7y4Ro3W7Mv5i2p81A/yG56oU1VYdNz9HS3KjndfbjTc7qA4DDrZ2PVJcnVPGO4RxJTf
sJcxgcH4HTyOvMCV6DGAODOcE42+Lmd0LU3CGYXeZfRcsS9PD3YX8tWFtiQdnSzTRMc6dVvsGTbo
RQKb6OC6Vco6NSBAwmHxmsNFnynu5u6zxFBZYlf6ir1amUlqq8HpEuQ5OQ4nbnQ6BYpjJyTodoVa
jttvPBiXrO0r8StcLzo0cC/2CCoA08vozD+otPkp3gc9ViaCvRAw3tMZ3DTUuKmgCQcx9ZYTD4/E
wUWXSVGc+N7knStXMKoHMfhMXXxSjaJ79d6KpqO3XIDJwrhtLdaue+T5+9qBceKR+s/8WmK1RgIt
5T8Trpry3rZ6jwG2iyUWYGLpHjU/W592hTkmv4FOT+cdki1Z4lb2FtlCzXhjpSInRz8cTEUbEXbu
6izfiKVXZyOAanwX3+Qqx4iqTlKbH8qJQ8cwkdXkzsyP3FPQ55jHZ0D2bTV2tfiR2IA015nAqjqO
BpqVP9sshkaO6AjJ2fG9Jepmc2JrLhabCNZlix0nZA+o7DqM6HivcRb5tdLxrpbjyogktmTZGOdF
BuzVhfHphU1sqac+UsgTIswAw15qKOgys/9b6cERHM4bPPVuuQ07ABU4jfbQ3YDDFwxkDmiic7sl
HDbvNgIzPtYN7zY9y2D/n14jGCgF4vVoQs8s/UvceYgd1KAyiTTCRhTomKWX50uY11PDUo2W2MI1
7FY/4z8jql1oOBrwMX0E0QVyB6vfpOkbB7pbpx54I8TuQfUBUKL1Dz4wHK7wtQhtPDzVTC4jGvVq
xN0XL5adxOeVrWguGsTAmwjnbAeuhqLrdtNmsP/oWO5hiBzfgxT9/Mttgi3+5UBkml0JYNId8H04
ELXLLbhwqA6btOL3uqz1K9AMXjj/xcYDuAulw7HuP04rFiz2UKgFeYagEzKHhBs2DGQ7IsHyNg5v
ftTfANrZgLTxd50HtOJAuWEiU37Y4AaQc9y1Con6+vkZXqqiLkK52S6CPfYm/NFJVli66EhKBxDX
E6IifhlhIttwsFhBKh/UFkTE/yGEFn5pqQpf6EJrwPp/U8PO7LHTBSPH+1RCHlMk2sCImVKU9+Nr
7LQNcSx6i+9N/RvjKD8TZeQTEg+38WyZFsNnj6rhTesYhxorjQdhhkRev9K9dK8haVbwPzrXZzGz
WY5qsQtHviG7VXGffX4rLMgfoGlrTGnQIXat0xne5wfLDqFuuW1h1nCj6nj+2cljss3RasNbrjaB
9znDXTHCYPdQ1FTtfWeUMAD6DMPez+NA9NLB/gfM5MipIuvjommwQAbMskLshYLePBixztHcFG2H
5k7VjmcA8J1r/vkfgJHk4HkBYT+xaGwv94umGVPZsrApmgyS1FJBr00SvZQV2Af+m/uyFnMtePIU
CdyCBx7fVoN82GQJV8YRx1cgd7w7QsmmHaZ8wjCYx5D0s+vhyr+1k5imaYZElJAS0Gbia5tlRK0z
oF2oHfbdpoN+s1QjKubPufNdAhmIjrfDZ37yZiv7H/LYn7BqN7L7RzkTT6tc4J0gzmJtg8I2LjXd
nttEwsYjAMOSeu+HoSUcof4laRtMSlfkEYh+/iZHSIntd0Ab5jvH4rhzefByHLNFNDz8nBJoWl8+
355LEGPOMz+NScu351BjGZKO/D2FNilxhqDFUU/YN4ER/Un+ita4+4/O3y6JN3Fo8h7zzO/YR0wn
1xEAWquU3LF+EKm7lI6p5h8WNZvXC4orBsAKpzH23zskSpiMOL6NtBClUp1ALjPMl602OsYvHLYi
Qs2umma4loiKaMqxqBZYBbLoOWPY9ObrEbUKzq2rnLqbaqid1WAevb8fUt9Pvn6vB2bKEzWIJz/Y
7VzdqmTI3PH+vYeFPiiLVaKYU+w3/lb5Sxoy05S4a73V7ayQZNwhjdaGmFKwl6+PuZyantGoXXb/
g4FS16tleY68PqElvngekQSVBGkWi1jtYpVICSALOOgW5jk0kZ6NlmQ0MVql1LuDJmBPMntcD2Ip
Kvng1rHabdjbHngx52AJzoMu8LUjxBV+NHMHuPJ9or6K1PBUKxI2LPyy8aKk0C/KRtZJdaPLUj/K
Uy1PKC1uGjk74fLIC+NABO+Jt4WfNSDZ9gH4PIjw1aEcODkB3s7mjnyyznqaPBtlEKEc/O3IeMYg
jyHODhTo6mrO2ohu5YtfGzNthrVcuAbufmSEFFHtiOzCUt8KBnVOY68jeoOi5sBKzslY4cLrtGY8
BqbhJq9N+tDPjsTiMMKU0LG4gRHN4nt6gg/KnG145x9JZUxQuBDDZIctEmgjS/oArD46zwcJVzX8
miqNCjf4R1OsJfwWiTGmmqNcBUh3IpTyYWPhXdV8T6uniq+7PKpbWnsIYVncB/+cpgBc8jqZsbOh
uMzf4vId05RNWKi88d72yeX1O0gWhX3kHLE96kc/MdMUpoQYdD220KEJcZvq5WzzQqYM5DZa3/bj
lwWHzaL4IzQESX5ZZleopAxQzEOzqMNi1gfB9aXvYKjKK6ZlWMBjr+Oe4glIz4AaccDPcbiwv33y
3Ufc3o5fFVLMF9y6e5c8BPT7VwkCFEgYT9YuC8SItn0A1viUZjePTQlVfb6lxK8i5hFuEJY6vlJ+
91llp1R/zfJrXFMBLfckOsKXflxEgqMFglne8cqbPyr8ajIQcx9E1LZ/fguE13YyrBeHAcbJoIDm
3dZBSQHW8nFeIgIo3E/HgSW8FW9BMWuoSsB09/9vYHkNw6aVmQ9z/Zb5UVDF3pPgfk11RBiJfPRQ
ajUex3KL0mFtYKnlBvHEGgvFA3S29dNVaRtS8sxg2xrv3ENBy+cK+2WvxFGXFzaEii8MhT2aR+m5
/gA0XTvNYInmvnolMqhuji/q4H21D0dGQpPymdi+rVitoJED3DFqqLfCHg1e5ju3/9Rfcz6kKs7B
3d9YgKMtFCpXPzXOIgTNF9lL9abBQK1I0wetdtp6tRPHFxmTXMVGRZUytYWg9/kLEdNp/X7wHPfI
OzMll2G19VhV45STbzuguW2BCl/hE8BvL/CreY8H7mpo2LgIBHtHUpB04q1iI7z7cG85ABqtGDUc
yNYQmeb1uae0fLMl+Ztq0Td4EiAj6GHZw/wESvDLb3opk6BGwTQB711yD0px6h4hgYJ9NvQwjlA7
+lbtoO3Jv1OfUyf8ziaUGtx1i8bswibWmHue0/BTJ6lDJApzYBuCA+V3JAgH1KgRV6Ckxk4UHnR6
HNlrsvyt/3fJJG4BKt/wkY0s98GHlsIrvY6WMBOjE2YRRwzUGcbwoUuxQdgg8q6+oXF9ND0b9TYI
WTfsyblmxeNdm/1PhbhcKvahgGUN1dvEJWgSfrK3/uEhVv0g63H7KcO+GcnWYm+hPTXqSSLMCVVS
dUbMVb4uP/y2U7zDBPFQDXSC639ng3mMv7jdcGi0OMCmPjryXFsRvbfqeCTDJDLXxQZzBRqbQA0y
CnJhjQEYqgdKoSBrpcdJ1HIrGJefvFqOZQvH590CjKbsvRqgAjqs5vA/TI17IfHaSKVXrUX70HtW
sutpMoKdNAsiWBo4JSNKXXUg+SViOvqySQVU9c7Ka2mWcQfr9ahqTa25yon1+3V9qCcDJFCkN6iL
8wZTg1X3FOXryKWI2rC20MSuwB0Le9LgPHNp3fudTaiYUuJfzMI65Y5w29SgpjVUJvyXhgrTyIKa
hLxPXvb//OrRnhoSrXr9emz/b9HOgyK+f2UIQCUIP/S5xIJnk5KW/ZWk7RIj2fXvKsHmAM2A0slj
nBDAnvXQK+t3uncfYmihQB2rMrI0rfkt9CWfKBYSptEsIfpDZmKyHfGwXz8blRqdtsQAQf2y+pZ5
NLhM2l4Kb2ND8hnL3ca6qmJEyEsLdJm5iKE4nS38moquaaWaINItKXQWLF7AzF2S7m6yoBC86JSg
qB4l+i4Xo39cv5cbzxa/7CahAmjjFYdIqGsy6EUW9DLhu9tT78zfQTjQ3GBSEph98ijth8q+gNLV
SqGiNyD2cVdEDJMbqY2M+WrTtc/FINNxQQQ1nn2TI87UATwvhBOWOVDBMkwSrmJn7B2HQo+oOPgr
SI20FNs3Atpk7kQsMA2VuH30CyvDqqEklV3jnfMATAcmzNegoHceJ3LPJ4OD0bIxJV8bxjQZLkjv
DwaugF0Z2l2dUcTNQ3ucoOzNQ1aLBRP22Q5sD56J5guT4v4EvE4wkKxq505M0xrOXmw6PjIXzyJb
qNm+eqRfeHpOdc2m4QKM5SM9IAf45JAdTl81RZKSkLQLqHq3oFoIvuyGUbWz4CHEX+BVjMvps4Tv
sKj2ZWD6c2eiIF5IFgox6OVL9t8wKe6jjA0nebkoQMB6rTvv9fXgVZxVnbLqvF+8QkJweA+x73Tt
TM0wlf0j5SNyolMm1EfOsjK+hkIRb8hpbwBANLuLYeIFLvXjVsZb7Et+L5Jf60aOnX+f6rVihmuf
sG0fwyeVsI0qOuBwAv3VPMuUt2sToQEm/L8IFFXehuEHtHo6RwTeZwZeY7MzSHrNOOGfYo/pFmsJ
DvvZGWi+Yk4DKGy8pyQtd9lisYQ/xobqyvEUgZij1RnKrGQQVsCkJ60JpBX82DYzOYKrERNVtxC5
sy6TKHiXwJCgy+JASmRGQz5HgP05EFfhVjpGaKUK1OwGCX3ug7wAJg4ogP0O3gnfwvBLEcTMCXsf
MC+aTGQxiIjHzEgfIw/IJzY+KvcmpY9pHTqeREy84OOQ6osdDtwPTiFwU0uf1hdGgeNI1HatXfaj
y8Of2PACMefekeV0rSNZ+XCUa+l0BWXSl2T2ht1ylMUp+VH8ipDM2cxyp28MUNxuWVY463mEr2WN
ijD9RjEqauBuBoeZH6RvxMILja672lwMP5z+PoWydBG8hJF/woLCcVlnmCcEZ2rq4zc3k5ThEQNH
ddgtjl1ItCs7HtgjYdnJixy2gEH8hk3FRATY8ZwFY3WfBzZT2xRadwPdvMOssH0ci3JB418jxduW
2GG71V3FDsW+i9smBEGtaKUC6+kxHDhFK7ndFdaLsaTdK12fNpQfDh6QH7Q2Vsw2I7/5Y6xcWXSc
P8liGRpRaFEIb9CzOvHgfbBPukBviGrNlXxFqsTD1L6F04oQByQI548qSHvnqhAKBnIfN+zQ9Tyo
ysZVpb/7na0+EKWUW1V5brlP3MvXHq6SyY/xB5eOjqvTShDeD2AKQu0UHCnoHH9PZDDYiL0uFSYc
4OXEHwUL4vD/fQw/4QimX1+I3kKHECg28dV4bV/q2bbIEy5SmKuxR8i+PbqYdJAOBPPe8uXL+0BS
OW/yIlzDSEnYkoAZn2qV33pwa/9AXQ8x77y8o1cqBAwLTtHwrIAvx6nI+DtWl2Nm1XYsOZ1pCDUe
kpCH9PnVqBwb0CtCptcDqF2GSyURiq0M/ExP2DYyLvsXDGjGLjXOafXhB26hx6nkyqO8kZnS8r3I
OIYiXF0Sm7z10AQfuXp2vk6Buvru2ShaaqF4SIUuwyUm0xOiLoXbXaJMROfLM4yTVzB/azEouywa
xDWitCoPxJzP6v6Hz1jfKoHbEsuBeFxCFnYtGRpUU9EXqSKIxlpCgKyCjrT75JzFvgmsyhtme++I
Xu1O4BX95ehsW6DigceI6Gi89jAG61pU34XT6KqdzAoV3g0tXsVQIsGKVHIUpRS+pvyNUB19PRnS
Ct8ftSqaBPOtxb7lCglZjbP1c1mlFunEkLhqYsUg4iFYRXhFUobCDzdAUIUc1eHVJCUjCStEZKPg
WJ5lkZWUh4PxLTrk5e7l1ttOr+6ayeRCIKTmRidt6/OfVDJyu4ZT9SO0nQGlWHCB6NghAcoswtPm
3lJaTSFrICdlFum+Xg6XbXn/Much8iSaqrYenrNQr3QzZtWp+P7PCpi0wacchZRvddK56L4y5t16
aXWWvCe57EdRWiF3mJOsL3ecycT5lAkvCiXxTDVd4v9Jx9adpaHBiOjTJixr+Okl+1aTSMr4mskF
vak2azZTXEcRBPcvx08ppLAWJkthqacVLdSV9aEDd47gbyhDE/ZsCxV8SgydNSle/yU+ZMBUACfz
9Y2Z+99kQdnZSSK2eDx4d2p6YSTCBwngDfK7HZwHeiHSU/RPvPQciDWFWBtF4uQFVRkPB+8gLArz
bY3EIwjnVq0GqLEFaxJO5IewdrCJmh+8/ClX2l4uj07oMlLDhgOAknRMIApql+O+ahXvovZju9ZS
yj2e3Ira9w5IwuZuxhvAgubE8k8QLWOqrm+39seL0O3xrF914pqxUJqmYRoi5MvQP3fPt6nPD4qa
xQrQhK6nyXKPam+mWLGPfQw8xmPunYWrPNqkrjwrPmqc19KsHTH1QwePXILT60s0LCuiW2A+RMQr
wtLZLfh5ZQWRE8eiDJrWAF2teM10yTCFYfiiAhmSxbedHnG+e9Ty2TNJ2qyRfDgs3m3JQJrGQ7un
luzj4bbM43y40ncdyGLBfu+mKU2UkL+g6HSR5Voi3s9LR7GcruzU0u3EAyXizOlMDC9gQ1EdMs72
rAXYNj+GufupY9S9XlkY1usBYEpI6/D6SubNnRBTfWIfS/Wto0SKYOGRbUgLOLNsEkWZtoyV4JIx
FkGZdPwu20eRY8pg4w7O/5QcwDwNJTRc6OoRlA9LQzfQq9Fl7hBpjfvu2Bq2HHeCxLH7DJ1cg2PQ
9WQceiwTj+7+r0ItdGoRLYhJAXco7xcXtIDobPSeraZ6Qgdttc2JIHO7Mz6cbwETMDDpBbqam+5G
+025zQn7eM+C29cR0RpivpMRqCgA+AUyTU/ouWiYmFjpI3fNFSAUQJfVVHeiEo5Tc8i6uwgA62eY
6DogzCTZ0vT3zej39hfccf/CkH+Flwz2mdElNOPTkXVHomFExV4Ye3VE6IBXb/57Bwl9GvEE+erI
d4tSi/zI5Ui0vyqcWY32VePO0xQC17meVG9Cl7X8vOY0rvlsw8kPLlPvQEzWQGx6GyOZC3NQvfn6
mTfJyUZuHpLZIcip0Kajr9qYr2sAmpaVm7RVAokxVmMzkmzhTt1Wsk+6uKJji/NmIYu8LJVHKsT7
Wp4ncb+cjgo8RK0VAY169mWREVRnqaybqMWm2i0FNB9luRVWEV7c5Qn5swRGPis2TK6SaOMn48ot
qcBTfbHs+/WqAkECEz+LakVDDRHUkszkub9oUaV17dAsAN0/+fXrMdaIU74DteDNmtTInXOcYA8i
amdPPnUvC/Y7opxsYERVX1eOw04gzge+TXgyQFosLEsphO2HMJRP2NUz79oQximh8iz2W+VNuVTF
88ck44twpgA9LED45EgjYGRrCkJ5ACp8/XwSjcwPGWmKCWTTOmaLBXKoUGFBPAQd33PQfptulWvd
/Iykkavp6zIa9CnFA7yOp/m7vyzCuZ8pRs6wq8LWZgJojzB7ABP7WnKe4SkiiHwYYu2akVIIZ/Zu
XjQuFUmzK/4oEUuvoY77+YLCMT1BhXCMPvPV1H4ZcmeRlGL4F5moreZ/s6eIsbMULTGuybQ2rDty
JAl6bOTOk+a3bhA1d+2VcN+YMJtTvmNW+CT0Ehyeppb2ek227gwCZz9iSrGsvFUQ8gfdMvenaI7K
YPzuyFIRdYZRO3mdUA2Muo+fUhuTMTcX7oaIQRVDZlszws9339V8mMzKTkp5z48JOmXx42la5aIl
f65NRtwDOL4EHOVYUL1MJh8TKvnMALPI4EG+8AXk2whgSJxT9mNs/0GeZf5w5GEr0LPJlriBztm1
d3DAVCd6D2BMb0gfoci6owu2LXH6pqGR0asGCio7FnJBQcpd+IG5KHazGK1FbqUIIi+T4qLP/PWS
IFVGdoC03nWHpwvxAWsE94Z1RnB3HNPrJmzSkq9P4CjZjhgmNQnVsSilYopzzlYVC9qYpWJdQVEh
lgSldho5I7R2IdL9lF9sl+DZ6/gzT1V3F0B/sny+U/kLRKZl2lLPDrwVBBWiy2H4Vmf1JPeBgh1q
4mGI8OAzZuLSEqvwHlb+nL4KL22JBsmXsIA9wqtbFX0MA8GThETQZmVyeQ9j8enceHz0+7hUaxqT
uMbuWW2UYiRjw6I9ToAkRfNVB8YcVP2T37zttxomCUrHo3IxDMqBsJpr5pYoe/J7j2s+0Se8yR8H
bBl7o/og01qZo3wF8AwcKLJjwPaIIALXKasRxR1WL2J7DOQ/nT5T6O/5OHIaWWimJOBMXWIZ5wUU
dD8etC6uav43veQE8yhtwG5w+GtMndEQxnFyQ/0NEzhhmZiUd1m81vKoE5qVEB1c0qr3VrY0zWsn
P6mtIx9i+9TSU3KW2beYqe4h/MFoEbdzqmOvfSEXPCbl0bpuMz0L20YClq5oNik8FtBrnlcH3YxU
5i1kcmEHmCyfvfwu9QF0q1NsNiTAQcPw/MF1k2cHZc99oEQICVyymSdJbla/NV7rbsCLkbIWnlP2
+qIU3/0E5yXGJaZ9n7XpyGOXUox09Pw+CrDcs+sb3NbxRBhDtW0NiXwy52Iq9dfLIfRcIbeYv6hL
/OaLnJfTWtwx9Q0yoDVAvGXS/biJTCKnjM0R3uyf4EN0vmKRkuJVKgmnwDG2Q1OqSB/oIGb/NYUE
RJVwYv7RX36e4zSSvacFSLiLEZDDDN1zWFSsKCTLxl0bZ1X+RU5NQioMQUBGufFZWX807fFHd1ed
qvyOmhgvoNT1CqUwrgWaSooTm9Zm3BSq+oSb7R3ioxctb/m2e93bcDT2qx5/CwzP3t9nKiWO51M+
ijH9AFL+Tab1kdmTjMx9gpefvk/MKMBPIA3jgZ/7wxL7zzBzLnCLcgSXkvnqj4V0C2JE1Eb2wmSN
N6AHaq6NzdCoTNQDQ/14xnnbFEnQ9Hsz5MpGZ7n+k3wTukhYPSSjByXT7npFKjhM/l9e4Jjl5I8J
YEuqH62gLHP/1XjTkCaRlzsg42oy1YFkYA+bP0qxUfjh0kQgSP/wkFU5vb0nUxLOYQk/gzfv1l9r
faogGNCQid0VuLJo629ZtDoodLD+gPNbxzhKtCPYSjRPQ+u8EY7CReZG5IVGzbTHm26W70B8vQEo
YTGJ6jGQVfKcfqoau8IGkZOaDqKzZvRCHsZ0LkwYE1JN9AqQLiVAma7fGvq2HjxtqAWCFlXQPGVI
SUGvoCvrs9XbM8pRK2SGlpRSVrfvNtCatsVMb76ZytAUJGyroa64O0KlCPdEsAPnqJdmhelMCR+D
dJYQVS4WooXPQBWWZjXxvEiWBAt01DOiB8wWyKOv9XD6ETnRXUtvv/CVQ30CvnMyhjj09dTV8v6s
dMJNzqjyfm/f/MMOJ1W6BkEOulIdxhpRbb7W8ax4My11LeKxppoILVwDy/kZuHE4CpUpP4pZ2YFD
Kmh9NpurSFwQNAdDiXxmC1Im0Xz5wNpjePgI3aIkXnFEd3YxsVWGNtzhXFk9TbDF0/t++tMkyzbm
kFP5Qqem+mzzod8FezUtrXXX2oFInL7F/F9ofkB+ZRFUNARPCbXbMLLYj0T1HN/0twrxNvvC1Tyv
vk70kAkwS3gfi3mDcOdpaKGxn4O4mi8WJ5RIzEi9kk0jRy3XRSotowqzhszfLDuL0iKluumc4GwE
hr9vSwvX14rxiiDAfiDyWYiDIrc29A116H1USkcPMdaPClowOtZDXwq8RLmdeHlC27K8v12gQV81
wPQa9HZZTa6k6duwRRtGMq8D5016RqY4aQNoVcUHNS8mbZlQWCnWQLCN2I1MXJMxN83qpVeQ6+Cf
U6utap+6D1uFQkFFycUPY1fclrQ3/3muO/khnANPwFmz0jVNv+cin7li/RGbRODilwA5/ezen1YT
R6KtXiCNAeGoIqpQZ7tED92MRB3XxdZ5axxzOJeAkrMMj5ZYyWtZTA39LcxlTB6T6dketBu49ttb
k5+n9Yj5iXUJkp9Rg5qi6QwmlfxECJHK7pqYi3SpDUNfPPo1zyOBwS3BHKssCV1cVKpE1r2+nI+S
H71gLOZ7I3+AHDiSJxQAtxLq4y4bM2M6lmNfk508qzNF9OucxXR5pv1C1iItX+vVaa0xvx55G0JA
556Q7fteTdygkytwliO8zMfLjSR3S6SSaKahoLklm942x2LILLXiwStSy8LzUiMkaP4uMgGmku90
r2kn2d8GJ6TzcBlk/YolpYQpZcCYnysdnDqZkIlOREF7bf0mxm7r5bFT9Jn9fx1T/tSXt5sUVm5n
ImCA8zkDAduRx7npQyGyuI1jYH+8EQpN9aVkc8k7KtakkpXcf7k5SkYGQLRdb4LqMiA0MYTS63Nm
UT4cS59KX6l4VX6Zd9CtdkyzgsVYleOrOfmwL1A44/JxOhdZXH9ZUSQOtTSwcg+SEL5xqQPgp72k
CntPHraUrr11H2tViwQhCaj2VKYFKQAOqM2ZNlP60Bx4IDlD3r941+UZHX5BYqhVxJdlQ/Iy3UQx
8o6SspMLZreLd5BIX5wQyQe1OvRuL77W6jPosJPsh10V1G7PfnibBE4sUdl08MeRBaGW42lvgUJh
pHkk4rv0AG6tGGBWdsUfzQ8n5NIKtj8E/+mJc1psnc2izxwu+5DidP8teMTUxppi0vvq8iMoXbMA
bYc+0y60tRQEuYE7pTP3eRlhC+GC7iOcqStPuRR8d7v6vUHPkJIdt9+0B7YSBRsV/Z4hp2ewKH3o
Vttb2gBXh8TIwiXWadW2ON3odjMK+zIPagmmNb+TbX5Nqsk9C3fbp20P8g8y+3FL5yyVm2W1sBvx
d1joE+zHrNQMCWKiW2dcs3ehet67DhJmO22bPkJ3WVQ8i7bi2yt310SLLVTsP2E1VyHvqoaagAGv
hUJuYAhTKDYdg6vkA7bCDLpVWk2kgU02yuF4c06VikOpbElJbaL/WDmmeAUkv3ogkseoBEyfqghT
hRa59XpYJMW10vPZLvZGRhD9Zz3CO9hnTTTP7SIKD/xW/Vyh2Kd3Kmg+p3cHD1/RaI9Fxqj0r5v4
inFdEHOQNBg8HwNqhkvNcrCRlXvfOJd+yz9yZAna
`pragma protect end_protected
