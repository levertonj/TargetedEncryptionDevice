// TEDv3_architecture.v

// Generated using ACDS version 14.1 190 at 2015.03.12.20:28:28

`timescale 1 ps / 1 ps
module TEDv3_architecture (
		output wire        black_interface_mac_mdio_connection_mdc,           //         black_interface_mac_mdio_connection.mdc
		input  wire        black_interface_mac_mdio_connection_mdio_in,       //                                            .mdio_in
		output wire        black_interface_mac_mdio_connection_mdio_out,      //                                            .mdio_out
		output wire        black_interface_mac_mdio_connection_mdio_oen,      //                                            .mdio_oen
		input  wire        black_interface_mac_misc_connection_xon_gen,       //         black_interface_mac_misc_connection.xon_gen
		input  wire        black_interface_mac_misc_connection_xoff_gen,      //                                            .xoff_gen
		input  wire        black_interface_mac_misc_connection_ff_tx_crc_fwd, //                                            .ff_tx_crc_fwd
		output wire        black_interface_mac_misc_connection_ff_tx_septy,   //                                            .ff_tx_septy
		output wire        black_interface_mac_misc_connection_tx_ff_uflow,   //                                            .tx_ff_uflow
		output wire        black_interface_mac_misc_connection_ff_tx_a_full,  //                                            .ff_tx_a_full
		output wire        black_interface_mac_misc_connection_ff_tx_a_empty, //                                            .ff_tx_a_empty
		output wire [17:0] black_interface_mac_misc_connection_rx_err_stat,   //                                            .rx_err_stat
		output wire [3:0]  black_interface_mac_misc_connection_rx_frm_type,   //                                            .rx_frm_type
		output wire        black_interface_mac_misc_connection_ff_rx_dsav,    //                                            .ff_rx_dsav
		output wire        black_interface_mac_misc_connection_ff_rx_a_full,  //                                            .ff_rx_a_full
		output wire        black_interface_mac_misc_connection_ff_rx_a_empty, //                                            .ff_rx_a_empty
		input  wire [3:0]  black_interface_mac_rgmii_connection_rgmii_in,     //        black_interface_mac_rgmii_connection.rgmii_in
		output wire [3:0]  black_interface_mac_rgmii_connection_rgmii_out,    //                                            .rgmii_out
		input  wire        black_interface_mac_rgmii_connection_rx_control,   //                                            .rx_control
		output wire        black_interface_mac_rgmii_connection_tx_control,   //                                            .tx_control
		input  wire        black_interface_mac_status_connection_set_10,      //       black_interface_mac_status_connection.set_10
		input  wire        black_interface_mac_status_connection_set_1000,    //                                            .set_1000
		output wire        black_interface_mac_status_connection_eth_mode,    //                                            .eth_mode
		output wire        black_interface_mac_status_connection_ena_10,      //                                            .ena_10
		input  wire        black_interface_pcs_mac_rx_clock_connection_clk,   // black_interface_pcs_mac_rx_clock_connection.clk
		input  wire        black_interface_pcs_mac_tx_clock_connection_clk,   // black_interface_pcs_mac_tx_clock_connection.clk
		input  wire        clk_clk,                                           //                                         clk.clk
		output wire [31:0] hex_conduit_hex_conduit,                           //                                 hex_conduit.hex_conduit
		input  wire [31:0] input_port_external_connection_export,             //              input_port_external_connection.export
		output wire [31:0] output_port_external_connection_export,            //             output_port_external_connection.export
		output wire        red_interface_mac_mdio_connection_mdc,             //           red_interface_mac_mdio_connection.mdc
		input  wire        red_interface_mac_mdio_connection_mdio_in,         //                                            .mdio_in
		output wire        red_interface_mac_mdio_connection_mdio_out,        //                                            .mdio_out
		output wire        red_interface_mac_mdio_connection_mdio_oen,        //                                            .mdio_oen
		input  wire        red_interface_mac_misc_connection_xon_gen,         //           red_interface_mac_misc_connection.xon_gen
		input  wire        red_interface_mac_misc_connection_xoff_gen,        //                                            .xoff_gen
		input  wire        red_interface_mac_misc_connection_ff_tx_crc_fwd,   //                                            .ff_tx_crc_fwd
		output wire        red_interface_mac_misc_connection_ff_tx_septy,     //                                            .ff_tx_septy
		output wire        red_interface_mac_misc_connection_tx_ff_uflow,     //                                            .tx_ff_uflow
		output wire        red_interface_mac_misc_connection_ff_tx_a_full,    //                                            .ff_tx_a_full
		output wire        red_interface_mac_misc_connection_ff_tx_a_empty,   //                                            .ff_tx_a_empty
		output wire [17:0] red_interface_mac_misc_connection_rx_err_stat,     //                                            .rx_err_stat
		output wire [3:0]  red_interface_mac_misc_connection_rx_frm_type,     //                                            .rx_frm_type
		output wire        red_interface_mac_misc_connection_ff_rx_dsav,      //                                            .ff_rx_dsav
		output wire        red_interface_mac_misc_connection_ff_rx_a_full,    //                                            .ff_rx_a_full
		output wire        red_interface_mac_misc_connection_ff_rx_a_empty,   //                                            .ff_rx_a_empty
		input  wire [3:0]  red_interface_mac_rgmii_connection_rgmii_in,       //          red_interface_mac_rgmii_connection.rgmii_in
		output wire [3:0]  red_interface_mac_rgmii_connection_rgmii_out,      //                                            .rgmii_out
		input  wire        red_interface_mac_rgmii_connection_rx_control,     //                                            .rx_control
		output wire        red_interface_mac_rgmii_connection_tx_control,     //                                            .tx_control
		input  wire        red_interface_mac_status_connection_set_10,        //         red_interface_mac_status_connection.set_10
		input  wire        red_interface_mac_status_connection_set_1000,      //                                            .set_1000
		output wire        red_interface_mac_status_connection_eth_mode,      //                                            .eth_mode
		output wire        red_interface_mac_status_connection_ena_10,        //                                            .ena_10
		input  wire        red_interface_pcs_mac_rx_clock_connection_clk,     //   red_interface_pcs_mac_rx_clock_connection.clk
		input  wire        red_interface_pcs_mac_tx_clock_connection_clk,     //   red_interface_pcs_mac_tx_clock_connection.clk
		input  wire        reset_reset_n                                      //                                       reset.reset_n
	);

	wire   [31:0] nios2_qsys_0_data_master_readdata;                                 // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire          nios2_qsys_0_data_master_waitrequest;                              // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire          nios2_qsys_0_data_master_debugaccess;                              // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [19:0] nios2_qsys_0_data_master_address;                                  // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire    [3:0] nios2_qsys_0_data_master_byteenable;                               // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire          nios2_qsys_0_data_master_read;                                     // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire          nios2_qsys_0_data_master_write;                                    // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire   [31:0] nios2_qsys_0_data_master_writedata;                                // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire   [31:0] red_interface_tx_mm_read_readdata;                                 // mm_interconnect_0:red_interface_tx_mm_read_readdata -> red_interface_tx:mm_read_readdata
	wire          red_interface_tx_mm_read_waitrequest;                              // mm_interconnect_0:red_interface_tx_mm_read_waitrequest -> red_interface_tx:mm_read_waitrequest
	wire   [31:0] red_interface_tx_mm_read_address;                                  // red_interface_tx:mm_read_address -> mm_interconnect_0:red_interface_tx_mm_read_address
	wire          red_interface_tx_mm_read_read;                                     // red_interface_tx:mm_read_read -> mm_interconnect_0:red_interface_tx_mm_read_read
	wire    [3:0] red_interface_tx_mm_read_byteenable;                               // red_interface_tx:mm_read_byteenable -> mm_interconnect_0:red_interface_tx_mm_read_byteenable
	wire          red_interface_tx_mm_read_readdatavalid;                            // mm_interconnect_0:red_interface_tx_mm_read_readdatavalid -> red_interface_tx:mm_read_readdatavalid
	wire    [4:0] red_interface_tx_mm_read_burstcount;                               // red_interface_tx:mm_read_burstcount -> mm_interconnect_0:red_interface_tx_mm_read_burstcount
	wire          black_interface_rx_mm_write_waitrequest;                           // mm_interconnect_0:black_interface_rx_mm_write_waitrequest -> black_interface_rx:mm_write_waitrequest
	wire   [31:0] black_interface_rx_mm_write_address;                               // black_interface_rx:mm_write_address -> mm_interconnect_0:black_interface_rx_mm_write_address
	wire    [3:0] black_interface_rx_mm_write_byteenable;                            // black_interface_rx:mm_write_byteenable -> mm_interconnect_0:black_interface_rx_mm_write_byteenable
	wire          black_interface_rx_mm_write_write;                                 // black_interface_rx:mm_write_write -> mm_interconnect_0:black_interface_rx_mm_write_write
	wire   [31:0] black_interface_rx_mm_write_writedata;                             // black_interface_rx:mm_write_writedata -> mm_interconnect_0:black_interface_rx_mm_write_writedata
	wire    [4:0] black_interface_rx_mm_write_burstcount;                            // black_interface_rx:mm_write_burstcount -> mm_interconnect_0:black_interface_rx_mm_write_burstcount
	wire   [31:0] ted_decryptor_read_master_readdata;                                // mm_interconnect_0:ted_decryptor_read_master_readdata -> ted_decryptor:avm_read_master_readdata
	wire          ted_decryptor_read_master_waitrequest;                             // mm_interconnect_0:ted_decryptor_read_master_waitrequest -> ted_decryptor:avm_read_master_waitrequest
	wire          ted_decryptor_read_master_read;                                    // ted_decryptor:avm_read_master_read -> mm_interconnect_0:ted_decryptor_read_master_read
	wire   [31:0] ted_decryptor_read_master_address;                                 // ted_decryptor:avm_read_master_address -> mm_interconnect_0:ted_decryptor_read_master_address
	wire          ted_decryptor_write_master_waitrequest;                            // mm_interconnect_0:ted_decryptor_write_master_waitrequest -> ted_decryptor:avm_write_master_waitrequest
	wire   [31:0] ted_decryptor_write_master_address;                                // ted_decryptor:avm_write_master_address -> mm_interconnect_0:ted_decryptor_write_master_address
	wire          ted_decryptor_write_master_write;                                  // ted_decryptor:avm_write_master_write -> mm_interconnect_0:ted_decryptor_write_master_write
	wire   [31:0] ted_decryptor_write_master_writedata;                              // ted_decryptor:avm_write_master_writedata -> mm_interconnect_0:ted_decryptor_write_master_writedata
	wire   [31:0] black_interface_tx_mm_read_readdata;                               // mm_interconnect_0:black_interface_tx_mm_read_readdata -> black_interface_tx:mm_read_readdata
	wire          black_interface_tx_mm_read_waitrequest;                            // mm_interconnect_0:black_interface_tx_mm_read_waitrequest -> black_interface_tx:mm_read_waitrequest
	wire   [31:0] black_interface_tx_mm_read_address;                                // black_interface_tx:mm_read_address -> mm_interconnect_0:black_interface_tx_mm_read_address
	wire          black_interface_tx_mm_read_read;                                   // black_interface_tx:mm_read_read -> mm_interconnect_0:black_interface_tx_mm_read_read
	wire    [3:0] black_interface_tx_mm_read_byteenable;                             // black_interface_tx:mm_read_byteenable -> mm_interconnect_0:black_interface_tx_mm_read_byteenable
	wire          black_interface_tx_mm_read_readdatavalid;                          // mm_interconnect_0:black_interface_tx_mm_read_readdatavalid -> black_interface_tx:mm_read_readdatavalid
	wire    [4:0] black_interface_tx_mm_read_burstcount;                             // black_interface_tx:mm_read_burstcount -> mm_interconnect_0:black_interface_tx_mm_read_burstcount
	wire          red_interface_rx_mm_write_waitrequest;                             // mm_interconnect_0:red_interface_rx_mm_write_waitrequest -> red_interface_rx:mm_write_waitrequest
	wire   [31:0] red_interface_rx_mm_write_address;                                 // red_interface_rx:mm_write_address -> mm_interconnect_0:red_interface_rx_mm_write_address
	wire    [3:0] red_interface_rx_mm_write_byteenable;                              // red_interface_rx:mm_write_byteenable -> mm_interconnect_0:red_interface_rx_mm_write_byteenable
	wire          red_interface_rx_mm_write_write;                                   // red_interface_rx:mm_write_write -> mm_interconnect_0:red_interface_rx_mm_write_write
	wire   [31:0] red_interface_rx_mm_write_writedata;                               // red_interface_rx:mm_write_writedata -> mm_interconnect_0:red_interface_rx_mm_write_writedata
	wire    [4:0] red_interface_rx_mm_write_burstcount;                              // red_interface_rx:mm_write_burstcount -> mm_interconnect_0:red_interface_rx_mm_write_burstcount
	wire   [31:0] ted_encryptor_read_master_readdata;                                // mm_interconnect_0:ted_encryptor_read_master_readdata -> ted_encryptor:avm_read_master_readdata
	wire          ted_encryptor_read_master_waitrequest;                             // mm_interconnect_0:ted_encryptor_read_master_waitrequest -> ted_encryptor:avm_read_master_waitrequest
	wire          ted_encryptor_read_master_read;                                    // ted_encryptor:avm_read_master_read -> mm_interconnect_0:ted_encryptor_read_master_read
	wire   [31:0] ted_encryptor_read_master_address;                                 // ted_encryptor:avm_read_master_address -> mm_interconnect_0:ted_encryptor_read_master_address
	wire          ted_encryptor_write_master_waitrequest;                            // mm_interconnect_0:ted_encryptor_write_master_waitrequest -> ted_encryptor:avm_write_master_waitrequest
	wire   [31:0] ted_encryptor_write_master_address;                                // ted_encryptor:avm_write_master_address -> mm_interconnect_0:ted_encryptor_write_master_address
	wire          ted_encryptor_write_master_write;                                  // ted_encryptor:avm_write_master_write -> mm_interconnect_0:ted_encryptor_write_master_write
	wire   [31:0] ted_encryptor_write_master_writedata;                              // ted_encryptor:avm_write_master_writedata -> mm_interconnect_0:ted_encryptor_write_master_writedata
	wire   [31:0] nios2_qsys_0_instruction_master_readdata;                          // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire          nios2_qsys_0_instruction_master_waitrequest;                       // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire   [19:0] nios2_qsys_0_instruction_master_address;                           // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire          nios2_qsys_0_instruction_master_read;                              // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire          mm_interconnect_0_hex_avalon_slave_0_chipselect;                   // mm_interconnect_0:hex_avalon_slave_0_chipselect -> hex:chipselect
	wire   [31:0] mm_interconnect_0_hex_avalon_slave_0_readdata;                     // hex:readdata -> mm_interconnect_0:hex_avalon_slave_0_readdata
	wire          mm_interconnect_0_hex_avalon_slave_0_read;                         // mm_interconnect_0:hex_avalon_slave_0_read -> hex:read
	wire    [3:0] mm_interconnect_0_hex_avalon_slave_0_byteenable;                   // mm_interconnect_0:hex_avalon_slave_0_byteenable -> hex:byteenable
	wire          mm_interconnect_0_hex_avalon_slave_0_write;                        // mm_interconnect_0:hex_avalon_slave_0_write -> hex:write
	wire   [31:0] mm_interconnect_0_hex_avalon_slave_0_writedata;                    // mm_interconnect_0:hex_avalon_slave_0_writedata -> hex:writedata
	wire   [31:0] mm_interconnect_0_black_interface_control_port_readdata;           // black_interface:reg_data_out -> mm_interconnect_0:black_interface_control_port_readdata
	wire          mm_interconnect_0_black_interface_control_port_waitrequest;        // black_interface:reg_busy -> mm_interconnect_0:black_interface_control_port_waitrequest
	wire    [7:0] mm_interconnect_0_black_interface_control_port_address;            // mm_interconnect_0:black_interface_control_port_address -> black_interface:reg_addr
	wire          mm_interconnect_0_black_interface_control_port_read;               // mm_interconnect_0:black_interface_control_port_read -> black_interface:reg_rd
	wire          mm_interconnect_0_black_interface_control_port_write;              // mm_interconnect_0:black_interface_control_port_write -> black_interface:reg_wr
	wire   [31:0] mm_interconnect_0_black_interface_control_port_writedata;          // mm_interconnect_0:black_interface_control_port_writedata -> black_interface:reg_data_in
	wire   [31:0] mm_interconnect_0_red_interface_control_port_readdata;             // red_interface:reg_data_out -> mm_interconnect_0:red_interface_control_port_readdata
	wire          mm_interconnect_0_red_interface_control_port_waitrequest;          // red_interface:reg_busy -> mm_interconnect_0:red_interface_control_port_waitrequest
	wire    [7:0] mm_interconnect_0_red_interface_control_port_address;              // mm_interconnect_0:red_interface_control_port_address -> red_interface:reg_addr
	wire          mm_interconnect_0_red_interface_control_port_read;                 // mm_interconnect_0:red_interface_control_port_read -> red_interface:reg_rd
	wire          mm_interconnect_0_red_interface_control_port_write;                // mm_interconnect_0:red_interface_control_port_write -> red_interface:reg_wr
	wire   [31:0] mm_interconnect_0_red_interface_control_port_writedata;            // mm_interconnect_0:red_interface_control_port_writedata -> red_interface:reg_data_in
	wire   [31:0] mm_interconnect_0_system_id_control_slave_readdata;                // system_id:readdata -> mm_interconnect_0:system_id_control_slave_readdata
	wire    [0:0] mm_interconnect_0_system_id_control_slave_address;                 // mm_interconnect_0:system_id_control_slave_address -> system_id:address
	wire   [31:0] mm_interconnect_0_ted_encryptor_csr_readdata;                      // ted_encryptor:avs_csr_readdata -> mm_interconnect_0:ted_encryptor_csr_readdata
	wire    [2:0] mm_interconnect_0_ted_encryptor_csr_address;                       // mm_interconnect_0:ted_encryptor_csr_address -> ted_encryptor:avs_csr_address
	wire          mm_interconnect_0_ted_encryptor_csr_write;                         // mm_interconnect_0:ted_encryptor_csr_write -> ted_encryptor:avs_csr_write
	wire   [31:0] mm_interconnect_0_ted_encryptor_csr_writedata;                     // mm_interconnect_0:ted_encryptor_csr_writedata -> ted_encryptor:avs_csr_writedata
	wire   [31:0] mm_interconnect_0_ted_decryptor_csr_readdata;                      // ted_decryptor:avs_csr_readdata -> mm_interconnect_0:ted_decryptor_csr_readdata
	wire    [2:0] mm_interconnect_0_ted_decryptor_csr_address;                       // mm_interconnect_0:ted_decryptor_csr_address -> ted_decryptor:avs_csr_address
	wire          mm_interconnect_0_ted_decryptor_csr_write;                         // mm_interconnect_0:ted_decryptor_csr_write -> ted_decryptor:avs_csr_write
	wire   [31:0] mm_interconnect_0_ted_decryptor_csr_writedata;                     // mm_interconnect_0:ted_decryptor_csr_writedata -> ted_decryptor:avs_csr_writedata
	wire   [31:0] mm_interconnect_0_red_interface_rx_csr_readdata;                   // red_interface_rx:csr_readdata -> mm_interconnect_0:red_interface_rx_csr_readdata
	wire    [2:0] mm_interconnect_0_red_interface_rx_csr_address;                    // mm_interconnect_0:red_interface_rx_csr_address -> red_interface_rx:csr_address
	wire          mm_interconnect_0_red_interface_rx_csr_read;                       // mm_interconnect_0:red_interface_rx_csr_read -> red_interface_rx:csr_read
	wire    [3:0] mm_interconnect_0_red_interface_rx_csr_byteenable;                 // mm_interconnect_0:red_interface_rx_csr_byteenable -> red_interface_rx:csr_byteenable
	wire          mm_interconnect_0_red_interface_rx_csr_write;                      // mm_interconnect_0:red_interface_rx_csr_write -> red_interface_rx:csr_write
	wire   [31:0] mm_interconnect_0_red_interface_rx_csr_writedata;                  // mm_interconnect_0:red_interface_rx_csr_writedata -> red_interface_rx:csr_writedata
	wire   [31:0] mm_interconnect_0_red_interface_tx_csr_readdata;                   // red_interface_tx:csr_readdata -> mm_interconnect_0:red_interface_tx_csr_readdata
	wire    [2:0] mm_interconnect_0_red_interface_tx_csr_address;                    // mm_interconnect_0:red_interface_tx_csr_address -> red_interface_tx:csr_address
	wire          mm_interconnect_0_red_interface_tx_csr_read;                       // mm_interconnect_0:red_interface_tx_csr_read -> red_interface_tx:csr_read
	wire    [3:0] mm_interconnect_0_red_interface_tx_csr_byteenable;                 // mm_interconnect_0:red_interface_tx_csr_byteenable -> red_interface_tx:csr_byteenable
	wire          mm_interconnect_0_red_interface_tx_csr_write;                      // mm_interconnect_0:red_interface_tx_csr_write -> red_interface_tx:csr_write
	wire   [31:0] mm_interconnect_0_red_interface_tx_csr_writedata;                  // mm_interconnect_0:red_interface_tx_csr_writedata -> red_interface_tx:csr_writedata
	wire   [31:0] mm_interconnect_0_black_interface_rx_csr_readdata;                 // black_interface_rx:csr_readdata -> mm_interconnect_0:black_interface_rx_csr_readdata
	wire    [2:0] mm_interconnect_0_black_interface_rx_csr_address;                  // mm_interconnect_0:black_interface_rx_csr_address -> black_interface_rx:csr_address
	wire          mm_interconnect_0_black_interface_rx_csr_read;                     // mm_interconnect_0:black_interface_rx_csr_read -> black_interface_rx:csr_read
	wire    [3:0] mm_interconnect_0_black_interface_rx_csr_byteenable;               // mm_interconnect_0:black_interface_rx_csr_byteenable -> black_interface_rx:csr_byteenable
	wire          mm_interconnect_0_black_interface_rx_csr_write;                    // mm_interconnect_0:black_interface_rx_csr_write -> black_interface_rx:csr_write
	wire   [31:0] mm_interconnect_0_black_interface_rx_csr_writedata;                // mm_interconnect_0:black_interface_rx_csr_writedata -> black_interface_rx:csr_writedata
	wire   [31:0] mm_interconnect_0_black_interface_tx_csr_readdata;                 // black_interface_tx:csr_readdata -> mm_interconnect_0:black_interface_tx_csr_readdata
	wire    [2:0] mm_interconnect_0_black_interface_tx_csr_address;                  // mm_interconnect_0:black_interface_tx_csr_address -> black_interface_tx:csr_address
	wire          mm_interconnect_0_black_interface_tx_csr_read;                     // mm_interconnect_0:black_interface_tx_csr_read -> black_interface_tx:csr_read
	wire    [3:0] mm_interconnect_0_black_interface_tx_csr_byteenable;               // mm_interconnect_0:black_interface_tx_csr_byteenable -> black_interface_tx:csr_byteenable
	wire          mm_interconnect_0_black_interface_tx_csr_write;                    // mm_interconnect_0:black_interface_tx_csr_write -> black_interface_tx:csr_write
	wire   [31:0] mm_interconnect_0_black_interface_tx_csr_writedata;                // mm_interconnect_0:black_interface_tx_csr_writedata -> black_interface_tx:csr_writedata
	wire          mm_interconnect_0_red_interface_rx_descriptor_slave_waitrequest;   // red_interface_rx:descriptor_slave_waitrequest -> mm_interconnect_0:red_interface_rx_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_red_interface_rx_descriptor_slave_byteenable;    // mm_interconnect_0:red_interface_rx_descriptor_slave_byteenable -> red_interface_rx:descriptor_slave_byteenable
	wire          mm_interconnect_0_red_interface_rx_descriptor_slave_write;         // mm_interconnect_0:red_interface_rx_descriptor_slave_write -> red_interface_rx:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_red_interface_rx_descriptor_slave_writedata;     // mm_interconnect_0:red_interface_rx_descriptor_slave_writedata -> red_interface_rx:descriptor_slave_writedata
	wire          mm_interconnect_0_red_interface_tx_descriptor_slave_waitrequest;   // red_interface_tx:descriptor_slave_waitrequest -> mm_interconnect_0:red_interface_tx_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_red_interface_tx_descriptor_slave_byteenable;    // mm_interconnect_0:red_interface_tx_descriptor_slave_byteenable -> red_interface_tx:descriptor_slave_byteenable
	wire          mm_interconnect_0_red_interface_tx_descriptor_slave_write;         // mm_interconnect_0:red_interface_tx_descriptor_slave_write -> red_interface_tx:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_red_interface_tx_descriptor_slave_writedata;     // mm_interconnect_0:red_interface_tx_descriptor_slave_writedata -> red_interface_tx:descriptor_slave_writedata
	wire          mm_interconnect_0_black_interface_rx_descriptor_slave_waitrequest; // black_interface_rx:descriptor_slave_waitrequest -> mm_interconnect_0:black_interface_rx_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_black_interface_rx_descriptor_slave_byteenable;  // mm_interconnect_0:black_interface_rx_descriptor_slave_byteenable -> black_interface_rx:descriptor_slave_byteenable
	wire          mm_interconnect_0_black_interface_rx_descriptor_slave_write;       // mm_interconnect_0:black_interface_rx_descriptor_slave_write -> black_interface_rx:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_black_interface_rx_descriptor_slave_writedata;   // mm_interconnect_0:black_interface_rx_descriptor_slave_writedata -> black_interface_rx:descriptor_slave_writedata
	wire          mm_interconnect_0_black_interface_tx_descriptor_slave_waitrequest; // black_interface_tx:descriptor_slave_waitrequest -> mm_interconnect_0:black_interface_tx_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_black_interface_tx_descriptor_slave_byteenable;  // mm_interconnect_0:black_interface_tx_descriptor_slave_byteenable -> black_interface_tx:descriptor_slave_byteenable
	wire          mm_interconnect_0_black_interface_tx_descriptor_slave_write;       // mm_interconnect_0:black_interface_tx_descriptor_slave_write -> black_interface_tx:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_black_interface_tx_descriptor_slave_writedata;   // mm_interconnect_0:black_interface_tx_descriptor_slave_writedata -> black_interface_tx:descriptor_slave_writedata
	wire   [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;         // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire          mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest;      // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire          mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess;      // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;          // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire          mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;             // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire    [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire          mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;            // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire   [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [31:0] mm_interconnect_0_red_interface_rx_response_readdata;              // red_interface_rx:response_readdata -> mm_interconnect_0:red_interface_rx_response_readdata
	wire          mm_interconnect_0_red_interface_rx_response_waitrequest;           // red_interface_rx:response_waitrequest -> mm_interconnect_0:red_interface_rx_response_waitrequest
	wire    [0:0] mm_interconnect_0_red_interface_rx_response_address;               // mm_interconnect_0:red_interface_rx_response_address -> red_interface_rx:response_address
	wire          mm_interconnect_0_red_interface_rx_response_read;                  // mm_interconnect_0:red_interface_rx_response_read -> red_interface_rx:response_read
	wire    [3:0] mm_interconnect_0_red_interface_rx_response_byteenable;            // mm_interconnect_0:red_interface_rx_response_byteenable -> red_interface_rx:response_byteenable
	wire   [31:0] mm_interconnect_0_black_interface_rx_response_readdata;            // black_interface_rx:response_readdata -> mm_interconnect_0:black_interface_rx_response_readdata
	wire          mm_interconnect_0_black_interface_rx_response_waitrequest;         // black_interface_rx:response_waitrequest -> mm_interconnect_0:black_interface_rx_response_waitrequest
	wire    [0:0] mm_interconnect_0_black_interface_rx_response_address;             // mm_interconnect_0:black_interface_rx_response_address -> black_interface_rx:response_address
	wire          mm_interconnect_0_black_interface_rx_response_read;                // mm_interconnect_0:black_interface_rx_response_read -> black_interface_rx:response_read
	wire    [3:0] mm_interconnect_0_black_interface_rx_response_byteenable;          // mm_interconnect_0:black_interface_rx_response_byteenable -> black_interface_rx:response_byteenable
	wire          mm_interconnect_0_output_port_s1_chipselect;                       // mm_interconnect_0:output_port_s1_chipselect -> output_port:chipselect
	wire   [31:0] mm_interconnect_0_output_port_s1_readdata;                         // output_port:readdata -> mm_interconnect_0:output_port_s1_readdata
	wire    [1:0] mm_interconnect_0_output_port_s1_address;                          // mm_interconnect_0:output_port_s1_address -> output_port:address
	wire          mm_interconnect_0_output_port_s1_write;                            // mm_interconnect_0:output_port_s1_write -> output_port:write_n
	wire   [31:0] mm_interconnect_0_output_port_s1_writedata;                        // mm_interconnect_0:output_port_s1_writedata -> output_port:writedata
	wire   [31:0] mm_interconnect_0_input_port_s1_readdata;                          // input_port:readdata -> mm_interconnect_0:input_port_s1_readdata
	wire    [1:0] mm_interconnect_0_input_port_s1_address;                           // mm_interconnect_0:input_port_s1_address -> input_port:address
	wire          mm_interconnect_0_instruction_memory_s1_chipselect;                // mm_interconnect_0:instruction_memory_s1_chipselect -> instruction_memory:chipselect
	wire   [31:0] mm_interconnect_0_instruction_memory_s1_readdata;                  // instruction_memory:readdata -> mm_interconnect_0:instruction_memory_s1_readdata
	wire   [15:0] mm_interconnect_0_instruction_memory_s1_address;                   // mm_interconnect_0:instruction_memory_s1_address -> instruction_memory:address
	wire    [3:0] mm_interconnect_0_instruction_memory_s1_byteenable;                // mm_interconnect_0:instruction_memory_s1_byteenable -> instruction_memory:byteenable
	wire          mm_interconnect_0_instruction_memory_s1_write;                     // mm_interconnect_0:instruction_memory_s1_write -> instruction_memory:write
	wire   [31:0] mm_interconnect_0_instruction_memory_s1_writedata;                 // mm_interconnect_0:instruction_memory_s1_writedata -> instruction_memory:writedata
	wire          mm_interconnect_0_instruction_memory_s1_clken;                     // mm_interconnect_0:instruction_memory_s1_clken -> instruction_memory:clken
	wire          mm_interconnect_0_heap_stack_s1_chipselect;                        // mm_interconnect_0:heap_stack_s1_chipselect -> heap_stack:chipselect
	wire   [31:0] mm_interconnect_0_heap_stack_s1_readdata;                          // heap_stack:readdata -> mm_interconnect_0:heap_stack_s1_readdata
	wire   [11:0] mm_interconnect_0_heap_stack_s1_address;                           // mm_interconnect_0:heap_stack_s1_address -> heap_stack:address
	wire    [3:0] mm_interconnect_0_heap_stack_s1_byteenable;                        // mm_interconnect_0:heap_stack_s1_byteenable -> heap_stack:byteenable
	wire          mm_interconnect_0_heap_stack_s1_write;                             // mm_interconnect_0:heap_stack_s1_write -> heap_stack:write
	wire   [31:0] mm_interconnect_0_heap_stack_s1_writedata;                         // mm_interconnect_0:heap_stack_s1_writedata -> heap_stack:writedata
	wire          mm_interconnect_0_heap_stack_s1_clken;                             // mm_interconnect_0:heap_stack_s1_clken -> heap_stack:clken
	wire          mm_interconnect_0_system_timer_s1_chipselect;                      // mm_interconnect_0:system_timer_s1_chipselect -> system_timer:chipselect
	wire   [15:0] mm_interconnect_0_system_timer_s1_readdata;                        // system_timer:readdata -> mm_interconnect_0:system_timer_s1_readdata
	wire    [3:0] mm_interconnect_0_system_timer_s1_address;                         // mm_interconnect_0:system_timer_s1_address -> system_timer:address
	wire          mm_interconnect_0_system_timer_s1_write;                           // mm_interconnect_0:system_timer_s1_write -> system_timer:write_n
	wire   [15:0] mm_interconnect_0_system_timer_s1_writedata;                       // mm_interconnect_0:system_timer_s1_writedata -> system_timer:writedata
	wire          mm_interconnect_0_performance_timer_s1_chipselect;                 // mm_interconnect_0:performance_timer_s1_chipselect -> performance_timer:chipselect
	wire   [15:0] mm_interconnect_0_performance_timer_s1_readdata;                   // performance_timer:readdata -> mm_interconnect_0:performance_timer_s1_readdata
	wire    [3:0] mm_interconnect_0_performance_timer_s1_address;                    // mm_interconnect_0:performance_timer_s1_address -> performance_timer:address
	wire          mm_interconnect_0_performance_timer_s1_write;                      // mm_interconnect_0:performance_timer_s1_write -> performance_timer:write_n
	wire   [15:0] mm_interconnect_0_performance_timer_s1_writedata;                  // mm_interconnect_0:performance_timer_s1_writedata -> performance_timer:writedata
	wire          mm_interconnect_0_red_to_black_memory_s1_chipselect;               // mm_interconnect_0:red_to_black_memory_s1_chipselect -> red_to_black_memory:chipselect
	wire   [31:0] mm_interconnect_0_red_to_black_memory_s1_readdata;                 // red_to_black_memory:readdata -> mm_interconnect_0:red_to_black_memory_s1_readdata
	wire   [12:0] mm_interconnect_0_red_to_black_memory_s1_address;                  // mm_interconnect_0:red_to_black_memory_s1_address -> red_to_black_memory:address
	wire    [3:0] mm_interconnect_0_red_to_black_memory_s1_byteenable;               // mm_interconnect_0:red_to_black_memory_s1_byteenable -> red_to_black_memory:byteenable
	wire          mm_interconnect_0_red_to_black_memory_s1_write;                    // mm_interconnect_0:red_to_black_memory_s1_write -> red_to_black_memory:write
	wire   [31:0] mm_interconnect_0_red_to_black_memory_s1_writedata;                // mm_interconnect_0:red_to_black_memory_s1_writedata -> red_to_black_memory:writedata
	wire          mm_interconnect_0_red_to_black_memory_s1_clken;                    // mm_interconnect_0:red_to_black_memory_s1_clken -> red_to_black_memory:clken
	wire          mm_interconnect_0_black_to_red_memory_s1_chipselect;               // mm_interconnect_0:black_to_red_memory_s1_chipselect -> black_to_red_memory:chipselect
	wire   [31:0] mm_interconnect_0_black_to_red_memory_s1_readdata;                 // black_to_red_memory:readdata -> mm_interconnect_0:black_to_red_memory_s1_readdata
	wire   [12:0] mm_interconnect_0_black_to_red_memory_s1_address;                  // mm_interconnect_0:black_to_red_memory_s1_address -> black_to_red_memory:address
	wire    [3:0] mm_interconnect_0_black_to_red_memory_s1_byteenable;               // mm_interconnect_0:black_to_red_memory_s1_byteenable -> black_to_red_memory:byteenable
	wire          mm_interconnect_0_black_to_red_memory_s1_write;                    // mm_interconnect_0:black_to_red_memory_s1_write -> black_to_red_memory:write
	wire   [31:0] mm_interconnect_0_black_to_red_memory_s1_writedata;                // mm_interconnect_0:black_to_red_memory_s1_writedata -> black_to_red_memory:writedata
	wire          mm_interconnect_0_black_to_red_memory_s1_clken;                    // mm_interconnect_0:black_to_red_memory_s1_clken -> black_to_red_memory:clken
	wire          irq_mapper_receiver0_irq;                                          // red_interface_rx:csr_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                          // red_interface_tx:csr_irq_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                          // black_interface_rx:csr_irq_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                          // black_interface_tx:csr_irq_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                          // system_timer:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                          // performance_timer:irq -> irq_mapper:receiver6_irq
	wire   [31:0] nios2_qsys_0_d_irq_irq;                                            // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire          red_interface_receive_valid;                                       // red_interface:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire   [31:0] red_interface_receive_data;                                        // red_interface:ff_rx_data -> avalon_st_adapter:in_0_data
	wire          red_interface_receive_ready;                                       // avalon_st_adapter:in_0_ready -> red_interface:ff_rx_rdy
	wire          red_interface_receive_startofpacket;                               // red_interface:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire          red_interface_receive_endofpacket;                                 // red_interface:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire    [5:0] red_interface_receive_error;                                       // red_interface:rx_err -> avalon_st_adapter:in_0_error
	wire    [1:0] red_interface_receive_empty;                                       // red_interface:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire          avalon_st_adapter_out_0_valid;                                     // avalon_st_adapter:out_0_valid -> red_interface_rx:st_sink_valid
	wire   [31:0] avalon_st_adapter_out_0_data;                                      // avalon_st_adapter:out_0_data -> red_interface_rx:st_sink_data
	wire          avalon_st_adapter_out_0_ready;                                     // red_interface_rx:st_sink_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                             // avalon_st_adapter:out_0_startofpacket -> red_interface_rx:st_sink_startofpacket
	wire          avalon_st_adapter_out_0_endofpacket;                               // avalon_st_adapter:out_0_endofpacket -> red_interface_rx:st_sink_endofpacket
	wire    [1:0] avalon_st_adapter_out_0_empty;                                     // avalon_st_adapter:out_0_empty -> red_interface_rx:st_sink_empty
	wire          black_interface_receive_valid;                                     // black_interface:ff_rx_dval -> avalon_st_adapter_001:in_0_valid
	wire   [31:0] black_interface_receive_data;                                      // black_interface:ff_rx_data -> avalon_st_adapter_001:in_0_data
	wire          black_interface_receive_ready;                                     // avalon_st_adapter_001:in_0_ready -> black_interface:ff_rx_rdy
	wire          black_interface_receive_startofpacket;                             // black_interface:ff_rx_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire          black_interface_receive_endofpacket;                               // black_interface:ff_rx_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire    [5:0] black_interface_receive_error;                                     // black_interface:rx_err -> avalon_st_adapter_001:in_0_error
	wire    [1:0] black_interface_receive_empty;                                     // black_interface:ff_rx_mod -> avalon_st_adapter_001:in_0_empty
	wire          avalon_st_adapter_001_out_0_valid;                                 // avalon_st_adapter_001:out_0_valid -> black_interface_rx:st_sink_valid
	wire   [31:0] avalon_st_adapter_001_out_0_data;                                  // avalon_st_adapter_001:out_0_data -> black_interface_rx:st_sink_data
	wire          avalon_st_adapter_001_out_0_ready;                                 // black_interface_rx:st_sink_ready -> avalon_st_adapter_001:out_0_ready
	wire          avalon_st_adapter_001_out_0_startofpacket;                         // avalon_st_adapter_001:out_0_startofpacket -> black_interface_rx:st_sink_startofpacket
	wire          avalon_st_adapter_001_out_0_endofpacket;                           // avalon_st_adapter_001:out_0_endofpacket -> black_interface_rx:st_sink_endofpacket
	wire    [1:0] avalon_st_adapter_001_out_0_empty;                                 // avalon_st_adapter_001:out_0_empty -> black_interface_rx:st_sink_empty
	wire          red_interface_tx_st_source_valid;                                  // red_interface_tx:st_source_valid -> avalon_st_adapter_002:in_0_valid
	wire   [31:0] red_interface_tx_st_source_data;                                   // red_interface_tx:st_source_data -> avalon_st_adapter_002:in_0_data
	wire          red_interface_tx_st_source_ready;                                  // avalon_st_adapter_002:in_0_ready -> red_interface_tx:st_source_ready
	wire          red_interface_tx_st_source_startofpacket;                          // red_interface_tx:st_source_startofpacket -> avalon_st_adapter_002:in_0_startofpacket
	wire          red_interface_tx_st_source_endofpacket;                            // red_interface_tx:st_source_endofpacket -> avalon_st_adapter_002:in_0_endofpacket
	wire    [1:0] red_interface_tx_st_source_empty;                                  // red_interface_tx:st_source_empty -> avalon_st_adapter_002:in_0_empty
	wire          avalon_st_adapter_002_out_0_valid;                                 // avalon_st_adapter_002:out_0_valid -> red_interface:ff_tx_wren
	wire   [31:0] avalon_st_adapter_002_out_0_data;                                  // avalon_st_adapter_002:out_0_data -> red_interface:ff_tx_data
	wire          avalon_st_adapter_002_out_0_ready;                                 // red_interface:ff_tx_rdy -> avalon_st_adapter_002:out_0_ready
	wire          avalon_st_adapter_002_out_0_startofpacket;                         // avalon_st_adapter_002:out_0_startofpacket -> red_interface:ff_tx_sop
	wire          avalon_st_adapter_002_out_0_endofpacket;                           // avalon_st_adapter_002:out_0_endofpacket -> red_interface:ff_tx_eop
	wire          avalon_st_adapter_002_out_0_error;                                 // avalon_st_adapter_002:out_0_error -> red_interface:ff_tx_err
	wire    [1:0] avalon_st_adapter_002_out_0_empty;                                 // avalon_st_adapter_002:out_0_empty -> red_interface:ff_tx_mod
	wire          black_interface_tx_st_source_valid;                                // black_interface_tx:st_source_valid -> avalon_st_adapter_003:in_0_valid
	wire   [31:0] black_interface_tx_st_source_data;                                 // black_interface_tx:st_source_data -> avalon_st_adapter_003:in_0_data
	wire          black_interface_tx_st_source_ready;                                // avalon_st_adapter_003:in_0_ready -> black_interface_tx:st_source_ready
	wire          black_interface_tx_st_source_startofpacket;                        // black_interface_tx:st_source_startofpacket -> avalon_st_adapter_003:in_0_startofpacket
	wire          black_interface_tx_st_source_endofpacket;                          // black_interface_tx:st_source_endofpacket -> avalon_st_adapter_003:in_0_endofpacket
	wire    [1:0] black_interface_tx_st_source_empty;                                // black_interface_tx:st_source_empty -> avalon_st_adapter_003:in_0_empty
	wire          avalon_st_adapter_003_out_0_valid;                                 // avalon_st_adapter_003:out_0_valid -> black_interface:ff_tx_wren
	wire   [31:0] avalon_st_adapter_003_out_0_data;                                  // avalon_st_adapter_003:out_0_data -> black_interface:ff_tx_data
	wire          avalon_st_adapter_003_out_0_ready;                                 // black_interface:ff_tx_rdy -> avalon_st_adapter_003:out_0_ready
	wire          avalon_st_adapter_003_out_0_startofpacket;                         // avalon_st_adapter_003:out_0_startofpacket -> black_interface:ff_tx_sop
	wire          avalon_st_adapter_003_out_0_endofpacket;                           // avalon_st_adapter_003:out_0_endofpacket -> black_interface:ff_tx_eop
	wire          avalon_st_adapter_003_out_0_error;                                 // avalon_st_adapter_003:out_0_error -> black_interface:ff_tx_err
	wire    [1:0] avalon_st_adapter_003_out_0_empty;                                 // avalon_st_adapter_003:out_0_empty -> black_interface:ff_tx_mod
	wire          rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, black_interface:reset, black_interface_rx:reset_n_reset_n, black_interface_tx:reset_n_reset_n, black_to_red_memory:reset, heap_stack:reset, hex:resetn, input_port:reset_n, instruction_memory:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, output_port:reset_n, performance_timer:reset_n, red_interface:reset, red_interface_rx:reset_n_reset_n, red_interface_tx:reset_n_reset_n, red_to_black_memory:reset, rst_translator:in_reset, system_id:reset_n, system_timer:reset_n, ted_decryptor:csi_clock_reset, ted_encryptor:csi_clock_reset]
	wire          rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [black_to_red_memory:reset_req, heap_stack:reset_req, instruction_memory:reset_req, nios2_qsys_0:reset_req, red_to_black_memory:reset_req, rst_translator:reset_req_in]
	wire          nios2_qsys_0_jtag_debug_module_reset_reset;                        // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	TEDv3_architecture_black_interface black_interface (
		.clk           (clk_clk),                                                    // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                             //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_black_interface_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_black_interface_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_black_interface_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_black_interface_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_black_interface_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_black_interface_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (black_interface_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (black_interface_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (black_interface_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (black_interface_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (black_interface_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (black_interface_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (black_interface_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (black_interface_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (black_interface_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (black_interface_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (clk_clk),                                                    //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                                    //     transmit_clock_connection.clk
		.ff_rx_data    (black_interface_receive_data),                               //                       receive.data
		.ff_rx_eop     (black_interface_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (black_interface_receive_error),                              //                              .error
		.ff_rx_mod     (black_interface_receive_empty),                              //                              .empty
		.ff_rx_rdy     (black_interface_receive_ready),                              //                              .ready
		.ff_rx_sop     (black_interface_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (black_interface_receive_valid),                              //                              .valid
		.ff_tx_data    (avalon_st_adapter_003_out_0_data),                           //                      transmit.data
		.ff_tx_eop     (avalon_st_adapter_003_out_0_endofpacket),                    //                              .endofpacket
		.ff_tx_err     (avalon_st_adapter_003_out_0_error),                          //                              .error
		.ff_tx_mod     (avalon_st_adapter_003_out_0_empty),                          //                              .empty
		.ff_tx_rdy     (avalon_st_adapter_003_out_0_ready),                          //                              .ready
		.ff_tx_sop     (avalon_st_adapter_003_out_0_startofpacket),                  //                              .startofpacket
		.ff_tx_wren    (avalon_st_adapter_003_out_0_valid),                          //                              .valid
		.mdc           (black_interface_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (black_interface_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (black_interface_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (black_interface_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.xon_gen       (black_interface_mac_misc_connection_xon_gen),                //           mac_misc_connection.xon_gen
		.xoff_gen      (black_interface_mac_misc_connection_xoff_gen),               //                              .xoff_gen
		.ff_tx_crc_fwd (black_interface_mac_misc_connection_ff_tx_crc_fwd),          //                              .ff_tx_crc_fwd
		.ff_tx_septy   (black_interface_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (black_interface_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (black_interface_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (black_interface_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (black_interface_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (black_interface_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (black_interface_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (black_interface_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (black_interface_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	TEDv3_architecture_black_interface_rx black_interface_rx (
		.clock_clk                    (clk_clk),                                                           //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                                   //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_black_interface_rx_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_black_interface_rx_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_black_interface_rx_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_black_interface_rx_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_black_interface_rx_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_black_interface_rx_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_black_interface_rx_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_black_interface_rx_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_black_interface_rx_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_black_interface_rx_descriptor_slave_byteenable),  //                 .byteenable
		.response_waitrequest         (mm_interconnect_0_black_interface_rx_response_waitrequest),         //         response.waitrequest
		.response_byteenable          (mm_interconnect_0_black_interface_rx_response_byteenable),          //                 .byteenable
		.response_address             (mm_interconnect_0_black_interface_rx_response_address),             //                 .address
		.response_readdata            (mm_interconnect_0_black_interface_rx_response_readdata),            //                 .readdata
		.response_read                (mm_interconnect_0_black_interface_rx_response_read),                //                 .read
		.csr_irq_irq                  (irq_mapper_receiver2_irq),                                          //          csr_irq.irq
		.mm_write_address             (black_interface_rx_mm_write_address),                               //         mm_write.address
		.mm_write_write               (black_interface_rx_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (black_interface_rx_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (black_interface_rx_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (black_interface_rx_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (black_interface_rx_mm_write_burstcount),                            //                 .burstcount
		.st_sink_data                 (avalon_st_adapter_001_out_0_data),                                  //          st_sink.data
		.st_sink_valid                (avalon_st_adapter_001_out_0_valid),                                 //                 .valid
		.st_sink_ready                (avalon_st_adapter_001_out_0_ready),                                 //                 .ready
		.st_sink_startofpacket        (avalon_st_adapter_001_out_0_startofpacket),                         //                 .startofpacket
		.st_sink_endofpacket          (avalon_st_adapter_001_out_0_endofpacket),                           //                 .endofpacket
		.st_sink_empty                (avalon_st_adapter_001_out_0_empty)                                  //                 .empty
	);

	TEDv3_architecture_black_interface_tx black_interface_tx (
		.clock_clk                    (clk_clk),                                                           //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                                   //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_black_interface_tx_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_black_interface_tx_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_black_interface_tx_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_black_interface_tx_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_black_interface_tx_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_black_interface_tx_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_black_interface_tx_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_black_interface_tx_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_black_interface_tx_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_black_interface_tx_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver3_irq),                                          //          csr_irq.irq
		.mm_read_address              (black_interface_tx_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (black_interface_tx_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (black_interface_tx_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (black_interface_tx_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (black_interface_tx_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (black_interface_tx_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (black_interface_tx_mm_read_burstcount),                             //                 .burstcount
		.st_source_data               (black_interface_tx_st_source_data),                                 //        st_source.data
		.st_source_valid              (black_interface_tx_st_source_valid),                                //                 .valid
		.st_source_ready              (black_interface_tx_st_source_ready),                                //                 .ready
		.st_source_startofpacket      (black_interface_tx_st_source_startofpacket),                        //                 .startofpacket
		.st_source_endofpacket        (black_interface_tx_st_source_endofpacket),                          //                 .endofpacket
		.st_source_empty              (black_interface_tx_st_source_empty)                                 //                 .empty
	);

	TEDv3_architecture_black_to_red_memory black_to_red_memory (
		.clk        (clk_clk),                                             //   clk1.clk
		.address    (mm_interconnect_0_black_to_red_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_black_to_red_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_black_to_red_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_black_to_red_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_black_to_red_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_black_to_red_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_black_to_red_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                   //       .reset_req
	);

	TEDv3_architecture_heap_stack heap_stack (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_heap_stack_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_heap_stack_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_heap_stack_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_heap_stack_s1_write),      //       .write
		.readdata   (mm_interconnect_0_heap_stack_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_heap_stack_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_heap_stack_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	reg32_avalon_interface hex (
		.read       (mm_interconnect_0_hex_avalon_slave_0_read),       // avalon_slave_0.read
		.write      (mm_interconnect_0_hex_avalon_slave_0_write),      //               .write
		.chipselect (mm_interconnect_0_hex_avalon_slave_0_chipselect), //               .chipselect
		.writedata  (mm_interconnect_0_hex_avalon_slave_0_writedata),  //               .writedata
		.byteenable (mm_interconnect_0_hex_avalon_slave_0_byteenable), //               .byteenable
		.readdata   (mm_interconnect_0_hex_avalon_slave_0_readdata),   //               .readdata
		.clock      (clk_clk),                                         //     clock_sink.clk
		.resetn     (~rst_controller_reset_out_reset),                 //     reset_sink.reset_n
		.Q_export   (hex_conduit_hex_conduit)                          //    conduit_end.hex_conduit
	);

	TEDv3_architecture_input_port input_port (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_input_port_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_input_port_s1_readdata), //                    .readdata
		.in_port  (input_port_external_connection_export)     // external_connection.export
	);

	TEDv3_architecture_instruction_memory instruction_memory (
		.clk        (clk_clk),                                            //   clk1.clk
		.address    (mm_interconnect_0_instruction_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_instruction_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_instruction_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_instruction_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_instruction_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_instruction_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_instruction_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                     // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                  //       .reset_req
	);

	TEDv3_architecture_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                   //               irq.irq
	);

	TEDv3_architecture_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	TEDv3_architecture_output_port output_port (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_output_port_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_output_port_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_output_port_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_output_port_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_output_port_s1_readdata),   //                    .readdata
		.out_port   (output_port_external_connection_export)       // external_connection.export
	);

	TEDv3_architecture_performance_timer performance_timer (
		.clk        (clk_clk),                                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   // reset.reset_n
		.address    (mm_interconnect_0_performance_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_performance_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_performance_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_performance_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_performance_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)                           //   irq.irq
	);

	TEDv3_architecture_black_interface red_interface (
		.clk           (clk_clk),                                                  // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                           //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_red_interface_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_red_interface_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_red_interface_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_red_interface_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_red_interface_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_red_interface_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (red_interface_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (red_interface_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (red_interface_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (red_interface_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (red_interface_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (red_interface_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (red_interface_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (red_interface_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (red_interface_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (red_interface_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (clk_clk),                                                  //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                                  //     transmit_clock_connection.clk
		.ff_rx_data    (red_interface_receive_data),                               //                       receive.data
		.ff_rx_eop     (red_interface_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (red_interface_receive_error),                              //                              .error
		.ff_rx_mod     (red_interface_receive_empty),                              //                              .empty
		.ff_rx_rdy     (red_interface_receive_ready),                              //                              .ready
		.ff_rx_sop     (red_interface_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (red_interface_receive_valid),                              //                              .valid
		.ff_tx_data    (avalon_st_adapter_002_out_0_data),                         //                      transmit.data
		.ff_tx_eop     (avalon_st_adapter_002_out_0_endofpacket),                  //                              .endofpacket
		.ff_tx_err     (avalon_st_adapter_002_out_0_error),                        //                              .error
		.ff_tx_mod     (avalon_st_adapter_002_out_0_empty),                        //                              .empty
		.ff_tx_rdy     (avalon_st_adapter_002_out_0_ready),                        //                              .ready
		.ff_tx_sop     (avalon_st_adapter_002_out_0_startofpacket),                //                              .startofpacket
		.ff_tx_wren    (avalon_st_adapter_002_out_0_valid),                        //                              .valid
		.mdc           (red_interface_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (red_interface_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (red_interface_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (red_interface_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.xon_gen       (red_interface_mac_misc_connection_xon_gen),                //           mac_misc_connection.xon_gen
		.xoff_gen      (red_interface_mac_misc_connection_xoff_gen),               //                              .xoff_gen
		.ff_tx_crc_fwd (red_interface_mac_misc_connection_ff_tx_crc_fwd),          //                              .ff_tx_crc_fwd
		.ff_tx_septy   (red_interface_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (red_interface_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (red_interface_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (red_interface_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (red_interface_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (red_interface_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (red_interface_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (red_interface_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (red_interface_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	TEDv3_architecture_red_interface_rx red_interface_rx (
		.clock_clk                    (clk_clk),                                                         //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                                 //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_red_interface_rx_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_red_interface_rx_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_red_interface_rx_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_red_interface_rx_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_red_interface_rx_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_red_interface_rx_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_red_interface_rx_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_red_interface_rx_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_red_interface_rx_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_red_interface_rx_descriptor_slave_byteenable),  //                 .byteenable
		.response_waitrequest         (mm_interconnect_0_red_interface_rx_response_waitrequest),         //         response.waitrequest
		.response_byteenable          (mm_interconnect_0_red_interface_rx_response_byteenable),          //                 .byteenable
		.response_address             (mm_interconnect_0_red_interface_rx_response_address),             //                 .address
		.response_readdata            (mm_interconnect_0_red_interface_rx_response_readdata),            //                 .readdata
		.response_read                (mm_interconnect_0_red_interface_rx_response_read),                //                 .read
		.csr_irq_irq                  (irq_mapper_receiver0_irq),                                        //          csr_irq.irq
		.mm_write_address             (red_interface_rx_mm_write_address),                               //         mm_write.address
		.mm_write_write               (red_interface_rx_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (red_interface_rx_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (red_interface_rx_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (red_interface_rx_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (red_interface_rx_mm_write_burstcount),                            //                 .burstcount
		.st_sink_data                 (avalon_st_adapter_out_0_data),                                    //          st_sink.data
		.st_sink_valid                (avalon_st_adapter_out_0_valid),                                   //                 .valid
		.st_sink_ready                (avalon_st_adapter_out_0_ready),                                   //                 .ready
		.st_sink_startofpacket        (avalon_st_adapter_out_0_startofpacket),                           //                 .startofpacket
		.st_sink_endofpacket          (avalon_st_adapter_out_0_endofpacket),                             //                 .endofpacket
		.st_sink_empty                (avalon_st_adapter_out_0_empty)                                    //                 .empty
	);

	TEDv3_architecture_black_interface_tx red_interface_tx (
		.clock_clk                    (clk_clk),                                                         //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                                 //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_red_interface_tx_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_red_interface_tx_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_red_interface_tx_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_red_interface_tx_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_red_interface_tx_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_red_interface_tx_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_red_interface_tx_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_red_interface_tx_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_red_interface_tx_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_red_interface_tx_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver1_irq),                                        //          csr_irq.irq
		.mm_read_address              (red_interface_tx_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (red_interface_tx_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (red_interface_tx_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (red_interface_tx_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (red_interface_tx_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (red_interface_tx_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (red_interface_tx_mm_read_burstcount),                             //                 .burstcount
		.st_source_data               (red_interface_tx_st_source_data),                                 //        st_source.data
		.st_source_valid              (red_interface_tx_st_source_valid),                                //                 .valid
		.st_source_ready              (red_interface_tx_st_source_ready),                                //                 .ready
		.st_source_startofpacket      (red_interface_tx_st_source_startofpacket),                        //                 .startofpacket
		.st_source_endofpacket        (red_interface_tx_st_source_endofpacket),                          //                 .endofpacket
		.st_source_empty              (red_interface_tx_st_source_empty)                                 //                 .empty
	);

	TEDv3_architecture_red_to_black_memory red_to_black_memory (
		.clk        (clk_clk),                                             //   clk1.clk
		.address    (mm_interconnect_0_red_to_black_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_red_to_black_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_red_to_black_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_red_to_black_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_red_to_black_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_red_to_black_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_red_to_black_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                   //       .reset_req
	);

	TEDv3_architecture_system_id system_id (
		.clock    (clk_clk),                                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //         reset.reset_n
		.readdata (mm_interconnect_0_system_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_system_id_control_slave_address)   //              .address
	);

	TEDv3_architecture_system_timer system_timer (
		.clk        (clk_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_system_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                      //   irq.irq
	);

	ted_crypto ted_decryptor (
		.csi_clock_clk                (clk_clk),                                       //        clock.clk
		.csi_clock_reset              (rst_controller_reset_out_reset),                //  clock_reset.reset
		.avm_read_master_read         (ted_decryptor_read_master_read),                //  read_master.read
		.avm_read_master_address      (ted_decryptor_read_master_address),             //             .address
		.avm_read_master_readdata     (ted_decryptor_read_master_readdata),            //             .readdata
		.avm_read_master_waitrequest  (ted_decryptor_read_master_waitrequest),         //             .waitrequest
		.avm_write_master_write       (ted_decryptor_write_master_write),              // write_master.write
		.avm_write_master_address     (ted_decryptor_write_master_address),            //             .address
		.avm_write_master_writedata   (ted_decryptor_write_master_writedata),          //             .writedata
		.avm_write_master_waitrequest (ted_decryptor_write_master_waitrequest),        //             .waitrequest
		.avs_csr_address              (mm_interconnect_0_ted_decryptor_csr_address),   //          csr.address
		.avs_csr_readdata             (mm_interconnect_0_ted_decryptor_csr_readdata),  //             .readdata
		.avs_csr_write                (mm_interconnect_0_ted_decryptor_csr_write),     //             .write
		.avs_csr_writedata            (mm_interconnect_0_ted_decryptor_csr_writedata)  //             .writedata
	);

	ted_crypto ted_encryptor (
		.csi_clock_clk                (clk_clk),                                       //        clock.clk
		.csi_clock_reset              (rst_controller_reset_out_reset),                //  clock_reset.reset
		.avm_read_master_read         (ted_encryptor_read_master_read),                //  read_master.read
		.avm_read_master_address      (ted_encryptor_read_master_address),             //             .address
		.avm_read_master_readdata     (ted_encryptor_read_master_readdata),            //             .readdata
		.avm_read_master_waitrequest  (ted_encryptor_read_master_waitrequest),         //             .waitrequest
		.avm_write_master_write       (ted_encryptor_write_master_write),              // write_master.write
		.avm_write_master_address     (ted_encryptor_write_master_address),            //             .address
		.avm_write_master_writedata   (ted_encryptor_write_master_writedata),          //             .writedata
		.avm_write_master_waitrequest (ted_encryptor_write_master_waitrequest),        //             .waitrequest
		.avs_csr_address              (mm_interconnect_0_ted_encryptor_csr_address),   //          csr.address
		.avs_csr_readdata             (mm_interconnect_0_ted_encryptor_csr_readdata),  //             .readdata
		.avs_csr_write                (mm_interconnect_0_ted_encryptor_csr_write),     //             .write
		.avs_csr_writedata            (mm_interconnect_0_ted_encryptor_csr_writedata)  //             .writedata
	);

	TEDv3_architecture_mm_interconnect_0 mm_interconnect_0 (
		.sys_clk_clk_clk                                  (clk_clk),                                                           //                                sys_clk_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                    // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.black_interface_rx_mm_write_address              (black_interface_rx_mm_write_address),                               //                black_interface_rx_mm_write.address
		.black_interface_rx_mm_write_waitrequest          (black_interface_rx_mm_write_waitrequest),                           //                                           .waitrequest
		.black_interface_rx_mm_write_burstcount           (black_interface_rx_mm_write_burstcount),                            //                                           .burstcount
		.black_interface_rx_mm_write_byteenable           (black_interface_rx_mm_write_byteenable),                            //                                           .byteenable
		.black_interface_rx_mm_write_write                (black_interface_rx_mm_write_write),                                 //                                           .write
		.black_interface_rx_mm_write_writedata            (black_interface_rx_mm_write_writedata),                             //                                           .writedata
		.black_interface_tx_mm_read_address               (black_interface_tx_mm_read_address),                                //                 black_interface_tx_mm_read.address
		.black_interface_tx_mm_read_waitrequest           (black_interface_tx_mm_read_waitrequest),                            //                                           .waitrequest
		.black_interface_tx_mm_read_burstcount            (black_interface_tx_mm_read_burstcount),                             //                                           .burstcount
		.black_interface_tx_mm_read_byteenable            (black_interface_tx_mm_read_byteenable),                             //                                           .byteenable
		.black_interface_tx_mm_read_read                  (black_interface_tx_mm_read_read),                                   //                                           .read
		.black_interface_tx_mm_read_readdata              (black_interface_tx_mm_read_readdata),                               //                                           .readdata
		.black_interface_tx_mm_read_readdatavalid         (black_interface_tx_mm_read_readdatavalid),                          //                                           .readdatavalid
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                                  //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                              //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                               //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                     //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                                 //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                                    //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                                //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                              //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                           //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                       //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                              //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                          //                                           .readdata
		.red_interface_rx_mm_write_address                (red_interface_rx_mm_write_address),                                 //                  red_interface_rx_mm_write.address
		.red_interface_rx_mm_write_waitrequest            (red_interface_rx_mm_write_waitrequest),                             //                                           .waitrequest
		.red_interface_rx_mm_write_burstcount             (red_interface_rx_mm_write_burstcount),                              //                                           .burstcount
		.red_interface_rx_mm_write_byteenable             (red_interface_rx_mm_write_byteenable),                              //                                           .byteenable
		.red_interface_rx_mm_write_write                  (red_interface_rx_mm_write_write),                                   //                                           .write
		.red_interface_rx_mm_write_writedata              (red_interface_rx_mm_write_writedata),                               //                                           .writedata
		.red_interface_tx_mm_read_address                 (red_interface_tx_mm_read_address),                                  //                   red_interface_tx_mm_read.address
		.red_interface_tx_mm_read_waitrequest             (red_interface_tx_mm_read_waitrequest),                              //                                           .waitrequest
		.red_interface_tx_mm_read_burstcount              (red_interface_tx_mm_read_burstcount),                               //                                           .burstcount
		.red_interface_tx_mm_read_byteenable              (red_interface_tx_mm_read_byteenable),                               //                                           .byteenable
		.red_interface_tx_mm_read_read                    (red_interface_tx_mm_read_read),                                     //                                           .read
		.red_interface_tx_mm_read_readdata                (red_interface_tx_mm_read_readdata),                                 //                                           .readdata
		.red_interface_tx_mm_read_readdatavalid           (red_interface_tx_mm_read_readdatavalid),                            //                                           .readdatavalid
		.ted_decryptor_read_master_address                (ted_decryptor_read_master_address),                                 //                  ted_decryptor_read_master.address
		.ted_decryptor_read_master_waitrequest            (ted_decryptor_read_master_waitrequest),                             //                                           .waitrequest
		.ted_decryptor_read_master_read                   (ted_decryptor_read_master_read),                                    //                                           .read
		.ted_decryptor_read_master_readdata               (ted_decryptor_read_master_readdata),                                //                                           .readdata
		.ted_decryptor_write_master_address               (ted_decryptor_write_master_address),                                //                 ted_decryptor_write_master.address
		.ted_decryptor_write_master_waitrequest           (ted_decryptor_write_master_waitrequest),                            //                                           .waitrequest
		.ted_decryptor_write_master_write                 (ted_decryptor_write_master_write),                                  //                                           .write
		.ted_decryptor_write_master_writedata             (ted_decryptor_write_master_writedata),                              //                                           .writedata
		.ted_encryptor_read_master_address                (ted_encryptor_read_master_address),                                 //                  ted_encryptor_read_master.address
		.ted_encryptor_read_master_waitrequest            (ted_encryptor_read_master_waitrequest),                             //                                           .waitrequest
		.ted_encryptor_read_master_read                   (ted_encryptor_read_master_read),                                    //                                           .read
		.ted_encryptor_read_master_readdata               (ted_encryptor_read_master_readdata),                                //                                           .readdata
		.ted_encryptor_write_master_address               (ted_encryptor_write_master_address),                                //                 ted_encryptor_write_master.address
		.ted_encryptor_write_master_waitrequest           (ted_encryptor_write_master_waitrequest),                            //                                           .waitrequest
		.ted_encryptor_write_master_write                 (ted_encryptor_write_master_write),                                  //                                           .write
		.ted_encryptor_write_master_writedata             (ted_encryptor_write_master_writedata),                              //                                           .writedata
		.black_interface_control_port_address             (mm_interconnect_0_black_interface_control_port_address),            //               black_interface_control_port.address
		.black_interface_control_port_write               (mm_interconnect_0_black_interface_control_port_write),              //                                           .write
		.black_interface_control_port_read                (mm_interconnect_0_black_interface_control_port_read),               //                                           .read
		.black_interface_control_port_readdata            (mm_interconnect_0_black_interface_control_port_readdata),           //                                           .readdata
		.black_interface_control_port_writedata           (mm_interconnect_0_black_interface_control_port_writedata),          //                                           .writedata
		.black_interface_control_port_waitrequest         (mm_interconnect_0_black_interface_control_port_waitrequest),        //                                           .waitrequest
		.black_interface_rx_csr_address                   (mm_interconnect_0_black_interface_rx_csr_address),                  //                     black_interface_rx_csr.address
		.black_interface_rx_csr_write                     (mm_interconnect_0_black_interface_rx_csr_write),                    //                                           .write
		.black_interface_rx_csr_read                      (mm_interconnect_0_black_interface_rx_csr_read),                     //                                           .read
		.black_interface_rx_csr_readdata                  (mm_interconnect_0_black_interface_rx_csr_readdata),                 //                                           .readdata
		.black_interface_rx_csr_writedata                 (mm_interconnect_0_black_interface_rx_csr_writedata),                //                                           .writedata
		.black_interface_rx_csr_byteenable                (mm_interconnect_0_black_interface_rx_csr_byteenable),               //                                           .byteenable
		.black_interface_rx_descriptor_slave_write        (mm_interconnect_0_black_interface_rx_descriptor_slave_write),       //        black_interface_rx_descriptor_slave.write
		.black_interface_rx_descriptor_slave_writedata    (mm_interconnect_0_black_interface_rx_descriptor_slave_writedata),   //                                           .writedata
		.black_interface_rx_descriptor_slave_byteenable   (mm_interconnect_0_black_interface_rx_descriptor_slave_byteenable),  //                                           .byteenable
		.black_interface_rx_descriptor_slave_waitrequest  (mm_interconnect_0_black_interface_rx_descriptor_slave_waitrequest), //                                           .waitrequest
		.black_interface_rx_response_address              (mm_interconnect_0_black_interface_rx_response_address),             //                black_interface_rx_response.address
		.black_interface_rx_response_read                 (mm_interconnect_0_black_interface_rx_response_read),                //                                           .read
		.black_interface_rx_response_readdata             (mm_interconnect_0_black_interface_rx_response_readdata),            //                                           .readdata
		.black_interface_rx_response_byteenable           (mm_interconnect_0_black_interface_rx_response_byteenable),          //                                           .byteenable
		.black_interface_rx_response_waitrequest          (mm_interconnect_0_black_interface_rx_response_waitrequest),         //                                           .waitrequest
		.black_interface_tx_csr_address                   (mm_interconnect_0_black_interface_tx_csr_address),                  //                     black_interface_tx_csr.address
		.black_interface_tx_csr_write                     (mm_interconnect_0_black_interface_tx_csr_write),                    //                                           .write
		.black_interface_tx_csr_read                      (mm_interconnect_0_black_interface_tx_csr_read),                     //                                           .read
		.black_interface_tx_csr_readdata                  (mm_interconnect_0_black_interface_tx_csr_readdata),                 //                                           .readdata
		.black_interface_tx_csr_writedata                 (mm_interconnect_0_black_interface_tx_csr_writedata),                //                                           .writedata
		.black_interface_tx_csr_byteenable                (mm_interconnect_0_black_interface_tx_csr_byteenable),               //                                           .byteenable
		.black_interface_tx_descriptor_slave_write        (mm_interconnect_0_black_interface_tx_descriptor_slave_write),       //        black_interface_tx_descriptor_slave.write
		.black_interface_tx_descriptor_slave_writedata    (mm_interconnect_0_black_interface_tx_descriptor_slave_writedata),   //                                           .writedata
		.black_interface_tx_descriptor_slave_byteenable   (mm_interconnect_0_black_interface_tx_descriptor_slave_byteenable),  //                                           .byteenable
		.black_interface_tx_descriptor_slave_waitrequest  (mm_interconnect_0_black_interface_tx_descriptor_slave_waitrequest), //                                           .waitrequest
		.black_to_red_memory_s1_address                   (mm_interconnect_0_black_to_red_memory_s1_address),                  //                     black_to_red_memory_s1.address
		.black_to_red_memory_s1_write                     (mm_interconnect_0_black_to_red_memory_s1_write),                    //                                           .write
		.black_to_red_memory_s1_readdata                  (mm_interconnect_0_black_to_red_memory_s1_readdata),                 //                                           .readdata
		.black_to_red_memory_s1_writedata                 (mm_interconnect_0_black_to_red_memory_s1_writedata),                //                                           .writedata
		.black_to_red_memory_s1_byteenable                (mm_interconnect_0_black_to_red_memory_s1_byteenable),               //                                           .byteenable
		.black_to_red_memory_s1_chipselect                (mm_interconnect_0_black_to_red_memory_s1_chipselect),               //                                           .chipselect
		.black_to_red_memory_s1_clken                     (mm_interconnect_0_black_to_red_memory_s1_clken),                    //                                           .clken
		.heap_stack_s1_address                            (mm_interconnect_0_heap_stack_s1_address),                           //                              heap_stack_s1.address
		.heap_stack_s1_write                              (mm_interconnect_0_heap_stack_s1_write),                             //                                           .write
		.heap_stack_s1_readdata                           (mm_interconnect_0_heap_stack_s1_readdata),                          //                                           .readdata
		.heap_stack_s1_writedata                          (mm_interconnect_0_heap_stack_s1_writedata),                         //                                           .writedata
		.heap_stack_s1_byteenable                         (mm_interconnect_0_heap_stack_s1_byteenable),                        //                                           .byteenable
		.heap_stack_s1_chipselect                         (mm_interconnect_0_heap_stack_s1_chipselect),                        //                                           .chipselect
		.heap_stack_s1_clken                              (mm_interconnect_0_heap_stack_s1_clken),                             //                                           .clken
		.hex_avalon_slave_0_write                         (mm_interconnect_0_hex_avalon_slave_0_write),                        //                         hex_avalon_slave_0.write
		.hex_avalon_slave_0_read                          (mm_interconnect_0_hex_avalon_slave_0_read),                         //                                           .read
		.hex_avalon_slave_0_readdata                      (mm_interconnect_0_hex_avalon_slave_0_readdata),                     //                                           .readdata
		.hex_avalon_slave_0_writedata                     (mm_interconnect_0_hex_avalon_slave_0_writedata),                    //                                           .writedata
		.hex_avalon_slave_0_byteenable                    (mm_interconnect_0_hex_avalon_slave_0_byteenable),                   //                                           .byteenable
		.hex_avalon_slave_0_chipselect                    (mm_interconnect_0_hex_avalon_slave_0_chipselect),                   //                                           .chipselect
		.input_port_s1_address                            (mm_interconnect_0_input_port_s1_address),                           //                              input_port_s1.address
		.input_port_s1_readdata                           (mm_interconnect_0_input_port_s1_readdata),                          //                                           .readdata
		.instruction_memory_s1_address                    (mm_interconnect_0_instruction_memory_s1_address),                   //                      instruction_memory_s1.address
		.instruction_memory_s1_write                      (mm_interconnect_0_instruction_memory_s1_write),                     //                                           .write
		.instruction_memory_s1_readdata                   (mm_interconnect_0_instruction_memory_s1_readdata),                  //                                           .readdata
		.instruction_memory_s1_writedata                  (mm_interconnect_0_instruction_memory_s1_writedata),                 //                                           .writedata
		.instruction_memory_s1_byteenable                 (mm_interconnect_0_instruction_memory_s1_byteenable),                //                                           .byteenable
		.instruction_memory_s1_chipselect                 (mm_interconnect_0_instruction_memory_s1_chipselect),                //                                           .chipselect
		.instruction_memory_s1_clken                      (mm_interconnect_0_instruction_memory_s1_clken),                     //                                           .clken
		.jtag_uart_avalon_jtag_slave_address              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),             //                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),               //                                           .write
		.jtag_uart_avalon_jtag_slave_read                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                //                                           .read
		.jtag_uart_avalon_jtag_slave_readdata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),            //                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),           //                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),         //                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),          //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),          //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),            //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),             //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),         //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),        //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),       //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest),      //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess),      //                                           .debugaccess
		.output_port_s1_address                           (mm_interconnect_0_output_port_s1_address),                          //                             output_port_s1.address
		.output_port_s1_write                             (mm_interconnect_0_output_port_s1_write),                            //                                           .write
		.output_port_s1_readdata                          (mm_interconnect_0_output_port_s1_readdata),                         //                                           .readdata
		.output_port_s1_writedata                         (mm_interconnect_0_output_port_s1_writedata),                        //                                           .writedata
		.output_port_s1_chipselect                        (mm_interconnect_0_output_port_s1_chipselect),                       //                                           .chipselect
		.performance_timer_s1_address                     (mm_interconnect_0_performance_timer_s1_address),                    //                       performance_timer_s1.address
		.performance_timer_s1_write                       (mm_interconnect_0_performance_timer_s1_write),                      //                                           .write
		.performance_timer_s1_readdata                    (mm_interconnect_0_performance_timer_s1_readdata),                   //                                           .readdata
		.performance_timer_s1_writedata                   (mm_interconnect_0_performance_timer_s1_writedata),                  //                                           .writedata
		.performance_timer_s1_chipselect                  (mm_interconnect_0_performance_timer_s1_chipselect),                 //                                           .chipselect
		.red_interface_control_port_address               (mm_interconnect_0_red_interface_control_port_address),              //                 red_interface_control_port.address
		.red_interface_control_port_write                 (mm_interconnect_0_red_interface_control_port_write),                //                                           .write
		.red_interface_control_port_read                  (mm_interconnect_0_red_interface_control_port_read),                 //                                           .read
		.red_interface_control_port_readdata              (mm_interconnect_0_red_interface_control_port_readdata),             //                                           .readdata
		.red_interface_control_port_writedata             (mm_interconnect_0_red_interface_control_port_writedata),            //                                           .writedata
		.red_interface_control_port_waitrequest           (mm_interconnect_0_red_interface_control_port_waitrequest),          //                                           .waitrequest
		.red_interface_rx_csr_address                     (mm_interconnect_0_red_interface_rx_csr_address),                    //                       red_interface_rx_csr.address
		.red_interface_rx_csr_write                       (mm_interconnect_0_red_interface_rx_csr_write),                      //                                           .write
		.red_interface_rx_csr_read                        (mm_interconnect_0_red_interface_rx_csr_read),                       //                                           .read
		.red_interface_rx_csr_readdata                    (mm_interconnect_0_red_interface_rx_csr_readdata),                   //                                           .readdata
		.red_interface_rx_csr_writedata                   (mm_interconnect_0_red_interface_rx_csr_writedata),                  //                                           .writedata
		.red_interface_rx_csr_byteenable                  (mm_interconnect_0_red_interface_rx_csr_byteenable),                 //                                           .byteenable
		.red_interface_rx_descriptor_slave_write          (mm_interconnect_0_red_interface_rx_descriptor_slave_write),         //          red_interface_rx_descriptor_slave.write
		.red_interface_rx_descriptor_slave_writedata      (mm_interconnect_0_red_interface_rx_descriptor_slave_writedata),     //                                           .writedata
		.red_interface_rx_descriptor_slave_byteenable     (mm_interconnect_0_red_interface_rx_descriptor_slave_byteenable),    //                                           .byteenable
		.red_interface_rx_descriptor_slave_waitrequest    (mm_interconnect_0_red_interface_rx_descriptor_slave_waitrequest),   //                                           .waitrequest
		.red_interface_rx_response_address                (mm_interconnect_0_red_interface_rx_response_address),               //                  red_interface_rx_response.address
		.red_interface_rx_response_read                   (mm_interconnect_0_red_interface_rx_response_read),                  //                                           .read
		.red_interface_rx_response_readdata               (mm_interconnect_0_red_interface_rx_response_readdata),              //                                           .readdata
		.red_interface_rx_response_byteenable             (mm_interconnect_0_red_interface_rx_response_byteenable),            //                                           .byteenable
		.red_interface_rx_response_waitrequest            (mm_interconnect_0_red_interface_rx_response_waitrequest),           //                                           .waitrequest
		.red_interface_tx_csr_address                     (mm_interconnect_0_red_interface_tx_csr_address),                    //                       red_interface_tx_csr.address
		.red_interface_tx_csr_write                       (mm_interconnect_0_red_interface_tx_csr_write),                      //                                           .write
		.red_interface_tx_csr_read                        (mm_interconnect_0_red_interface_tx_csr_read),                       //                                           .read
		.red_interface_tx_csr_readdata                    (mm_interconnect_0_red_interface_tx_csr_readdata),                   //                                           .readdata
		.red_interface_tx_csr_writedata                   (mm_interconnect_0_red_interface_tx_csr_writedata),                  //                                           .writedata
		.red_interface_tx_csr_byteenable                  (mm_interconnect_0_red_interface_tx_csr_byteenable),                 //                                           .byteenable
		.red_interface_tx_descriptor_slave_write          (mm_interconnect_0_red_interface_tx_descriptor_slave_write),         //          red_interface_tx_descriptor_slave.write
		.red_interface_tx_descriptor_slave_writedata      (mm_interconnect_0_red_interface_tx_descriptor_slave_writedata),     //                                           .writedata
		.red_interface_tx_descriptor_slave_byteenable     (mm_interconnect_0_red_interface_tx_descriptor_slave_byteenable),    //                                           .byteenable
		.red_interface_tx_descriptor_slave_waitrequest    (mm_interconnect_0_red_interface_tx_descriptor_slave_waitrequest),   //                                           .waitrequest
		.red_to_black_memory_s1_address                   (mm_interconnect_0_red_to_black_memory_s1_address),                  //                     red_to_black_memory_s1.address
		.red_to_black_memory_s1_write                     (mm_interconnect_0_red_to_black_memory_s1_write),                    //                                           .write
		.red_to_black_memory_s1_readdata                  (mm_interconnect_0_red_to_black_memory_s1_readdata),                 //                                           .readdata
		.red_to_black_memory_s1_writedata                 (mm_interconnect_0_red_to_black_memory_s1_writedata),                //                                           .writedata
		.red_to_black_memory_s1_byteenable                (mm_interconnect_0_red_to_black_memory_s1_byteenable),               //                                           .byteenable
		.red_to_black_memory_s1_chipselect                (mm_interconnect_0_red_to_black_memory_s1_chipselect),               //                                           .chipselect
		.red_to_black_memory_s1_clken                     (mm_interconnect_0_red_to_black_memory_s1_clken),                    //                                           .clken
		.system_id_control_slave_address                  (mm_interconnect_0_system_id_control_slave_address),                 //                    system_id_control_slave.address
		.system_id_control_slave_readdata                 (mm_interconnect_0_system_id_control_slave_readdata),                //                                           .readdata
		.system_timer_s1_address                          (mm_interconnect_0_system_timer_s1_address),                         //                            system_timer_s1.address
		.system_timer_s1_write                            (mm_interconnect_0_system_timer_s1_write),                           //                                           .write
		.system_timer_s1_readdata                         (mm_interconnect_0_system_timer_s1_readdata),                        //                                           .readdata
		.system_timer_s1_writedata                        (mm_interconnect_0_system_timer_s1_writedata),                       //                                           .writedata
		.system_timer_s1_chipselect                       (mm_interconnect_0_system_timer_s1_chipselect),                      //                                           .chipselect
		.ted_decryptor_csr_address                        (mm_interconnect_0_ted_decryptor_csr_address),                       //                          ted_decryptor_csr.address
		.ted_decryptor_csr_write                          (mm_interconnect_0_ted_decryptor_csr_write),                         //                                           .write
		.ted_decryptor_csr_readdata                       (mm_interconnect_0_ted_decryptor_csr_readdata),                      //                                           .readdata
		.ted_decryptor_csr_writedata                      (mm_interconnect_0_ted_decryptor_csr_writedata),                     //                                           .writedata
		.ted_encryptor_csr_address                        (mm_interconnect_0_ted_encryptor_csr_address),                       //                          ted_encryptor_csr.address
		.ted_encryptor_csr_write                          (mm_interconnect_0_ted_encryptor_csr_write),                         //                                           .write
		.ted_encryptor_csr_readdata                       (mm_interconnect_0_ted_encryptor_csr_readdata),                      //                                           .readdata
		.ted_encryptor_csr_writedata                      (mm_interconnect_0_ted_encryptor_csr_writedata)                      //                                           .writedata
	);

	TEDv3_architecture_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	TEDv3_architecture_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (red_interface_receive_data),            //     in_0.data
		.in_0_valid          (red_interface_receive_valid),           //         .valid
		.in_0_ready          (red_interface_receive_ready),           //         .ready
		.in_0_startofpacket  (red_interface_receive_startofpacket),   //         .startofpacket
		.in_0_endofpacket    (red_interface_receive_endofpacket),     //         .endofpacket
		.in_0_empty          (red_interface_receive_empty),           //         .empty
		.in_0_error          (red_interface_receive_error),           //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)          //         .empty
	);

	TEDv3_architecture_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (black_interface_receive_data),              //     in_0.data
		.in_0_valid          (black_interface_receive_valid),             //         .valid
		.in_0_ready          (black_interface_receive_ready),             //         .ready
		.in_0_startofpacket  (black_interface_receive_startofpacket),     //         .startofpacket
		.in_0_endofpacket    (black_interface_receive_endofpacket),       //         .endofpacket
		.in_0_empty          (black_interface_receive_empty),             //         .empty
		.in_0_error          (black_interface_receive_error),             //         .error
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)          //         .empty
	);

	TEDv3_architecture_avalon_st_adapter_002 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_002 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (red_interface_tx_st_source_data),           //     in_0.data
		.in_0_valid          (red_interface_tx_st_source_valid),          //         .valid
		.in_0_ready          (red_interface_tx_st_source_ready),          //         .ready
		.in_0_startofpacket  (red_interface_tx_st_source_startofpacket),  //         .startofpacket
		.in_0_endofpacket    (red_interface_tx_st_source_endofpacket),    //         .endofpacket
		.in_0_empty          (red_interface_tx_st_source_empty),          //         .empty
		.out_0_data          (avalon_st_adapter_002_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_002_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_002_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_002_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_002_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_002_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_002_out_0_error)          //         .error
	);

	TEDv3_architecture_avalon_st_adapter_002 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_003 (
		.in_clk_0_clk        (clk_clk),                                    // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),             // in_rst_0.reset
		.in_0_data           (black_interface_tx_st_source_data),          //     in_0.data
		.in_0_valid          (black_interface_tx_st_source_valid),         //         .valid
		.in_0_ready          (black_interface_tx_st_source_ready),         //         .ready
		.in_0_startofpacket  (black_interface_tx_st_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (black_interface_tx_st_source_endofpacket),   //         .endofpacket
		.in_0_empty          (black_interface_tx_st_source_empty),         //         .empty
		.out_0_data          (avalon_st_adapter_003_out_0_data),           //    out_0.data
		.out_0_valid         (avalon_st_adapter_003_out_0_valid),          //         .valid
		.out_0_ready         (avalon_st_adapter_003_out_0_ready),          //         .ready
		.out_0_startofpacket (avalon_st_adapter_003_out_0_startofpacket),  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_003_out_0_endofpacket),    //         .endofpacket
		.out_0_empty         (avalon_st_adapter_003_out_0_empty),          //         .empty
		.out_0_error         (avalon_st_adapter_003_out_0_error)           //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
